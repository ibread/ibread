//# 3 inputs
//# 6 outputs
//# 14 D-type flipflops
//# 44 inverters
//# 75 gates (31 ANDs + 9 NANDs + 16 ORs + 19 NORs)

module dff (CK,Q,D);
input CK,D;
output Q;

  wire NM,NCK;
  trireg NQ,M;

  nmos N7 (M,D,NCK);
  not P3 (NM,M);
  nmos N9 (NQ,NM,CK);
  not P5 (Q,NQ);
  not P1 (NCK,CK);

endmodule

module s298 (scan_enable, scan_data_in, send_CK, send_GND, send_VDD, recv_CK, recv_GND, recv_VDD, hsend_G0, hsend_G1, hsend_G2, scan_data_out, hrecv_G117, hrecv_G132, hrecv_G66, hrecv_G118, hrecv_G133, hrecv_G67, hsend_G118, hsend_G133, hsend_G67);

input scan_enable, scan_data_in, send_CK, send_GND, send_VDD, recv_CK, recv_GND, recv_VDD, hsend_G0, hsend_G1, hsend_G2;

wire send_G0, send_G1, send_G2, recv_G0, recv_G1, recv_G2, send_G117, send_G132, send_G66, send_G118, send_G133, send_G67, recv_G117, recv_G132, recv_G66, recv_G118, recv_G133, recv_G67, send_G10, send_G29, send_G11, send_G30, send_G12, send_G34, send_G13, send_G39, send_G14, send_G44, send_G15, send_G56, send_G16, send_G86, send_G17, send_G92, send_G18, send_G98, send_G19, send_G102, send_G20, send_G107, send_G21, send_G113, send_G22, send_G119, send_G23, send_G125, send_G28, send_G130, send_G38, send_G40, send_G45, send_G46, send_G50, send_G51, send_G54, send_G55, send_G59, send_G60, send_G64, send_II155, send_II158, send_G76, send_G82, send_G87, send_G91, send_G93, send_G96, send_G99, send_G103, send_G108, send_G112, send_G114, send_II210, send_II213, send_G120, send_G124, send_G121, send_II221, send_G126, send_G131, send_G127, send_II229, send_II232, send_II235, send_II238, send_G26, send_G27, send_G31, send_G32, send_G33, send_G35, send_G36, send_G37, send_G42, send_G41, send_G48, send_G47, send_G49, send_G52, send_G57, send_G61, send_G58, send_G65, send_G62, send_G63, send_G74, send_G75, send_G88, send_G89, send_G90, send_G94, send_G95, send_G100, send_G105, send_G104, send_G110, send_G109, send_G111, send_G115, send_G122, send_G123, send_G128, send_G129, send_G24, send_G25, send_G68, send_G69, send_G70, send_G71, send_G72, send_G73, send_G77, send_G78, send_G79, send_G80, send_G81, send_G83, send_G84, send_G85, send_G43, send_G97, send_G101, send_G106, send_G116, send_G53, recv_G10, recv_G29, recv_G11, recv_G30, recv_G12, recv_G34, recv_G13, recv_G39, recv_G14, recv_G44, recv_G15, recv_G56, recv_G16, recv_G86, recv_G17, recv_G92, recv_G18, recv_G98, recv_G19, recv_G102, recv_G20, recv_G107, recv_G21, recv_G113, recv_G22, recv_G119, recv_G23, recv_G125, recv_G28, recv_G130, recv_G38, recv_G40, recv_G45, recv_G46, recv_G50, recv_G51, recv_G54, recv_G55, recv_G59, recv_G60, recv_G64, recv_II155, recv_II158, recv_G76, recv_G82, recv_G87, recv_G91, recv_G93, recv_G96, recv_G99, recv_G103, recv_G108, recv_G112, recv_G114, recv_II210, recv_II213, recv_G120, recv_G124, recv_G121, recv_II221, recv_G126, recv_G131, recv_G127, recv_II229, recv_II232, recv_II235, recv_II238, recv_G26, recv_G27, recv_G31, recv_G32, recv_G33, recv_G35, recv_G36, recv_G37, recv_G42, recv_G41, recv_G48, recv_G47, recv_G49, recv_G52, recv_G57, recv_G61, recv_G58, recv_G65, recv_G62, recv_G63, recv_G74, recv_G75, recv_G88, recv_G89, recv_G90, recv_G94, recv_G95, recv_G100, recv_G105, recv_G104, recv_G110, recv_G109, recv_G111, recv_G115, recv_G122, recv_G123, recv_G128, recv_G129, recv_G24, recv_G25, recv_G68, recv_G69, recv_G70, recv_G71, recv_G72, recv_G73, recv_G77, recv_G78, recv_G79, recv_G80, recv_G81, recv_G83, recv_G84, recv_G85, recv_G43, recv_G97, recv_G101, recv_G106, recv_G116, recv_G53;

output scan_data_out, hrecv_G117, hrecv_G132, hrecv_G66, hrecv_G118, hrecv_G133, hrecv_G67, hsend_G118, hsend_G133, hsend_G67;


// scan chain begins here

SDFFNSR MID_DFF0(.CK(send_CK), .D(SEND_G117), .Q(RECV_HG0), .SI(scan_data_in), .SE(scan_enable));
SDFFNSR MID_DFF1(.CK(send_CK), .D(SEND_G132), .Q(RECV_HG1), .SI(RECV_HG0), .SE(scan_enable));
SDFFNSR MID_DFF2(.CK(send_CK), .D(SEND_G66), .Q(RECV_HG2), .SI(RECV_HG1), .SE(scan_enable));
SDFFNSR SEND_I_DFF0(.CK(send_CK), .D(hsend_G0), .Q(send_G0), .SI(RECV_HG2), .SE(scan_enable));
SDFFNSR SEND_I_DFF1(.CK(send_CK), .D(hsend_G1), .Q(send_G1), .SI(send_G0), .SE(scan_enable));
SDFFNSR SEND_I_DFF2(.CK(send_CK), .D(hsend_G2), .Q(send_G2), .SI(send_G1), .SE(scan_enable));
SDFFNSR SEND_O_DFF3(.CK(send_CK), .D(send_G118), .Q(hsend_G118), .SI(send_G2), .SE(scan_enable));
SDFFNSR SEND_O_DFF4(.CK(send_CK), .D(send_G133), .Q(hsend_G133), .SI(hsend_G118), .SE(scan_enable));
SDFFNSR SEND_O_DFF5(.CK(send_CK), .D(send_G67), .Q(hsend_G67), .SI(hsend_G133), .SE(scan_enable));
SDFFNSR RECV_I_DFF0(.CK(recv_CK), .D(hrecv_G0), .Q(recv_G0), .SI(hsend_G67), .SE(scan_enable));
SDFFNSR RECV_I_DFF1(.CK(recv_CK), .D(hrecv_G1), .Q(recv_G1), .SI(recv_G0), .SE(scan_enable));
SDFFNSR RECV_I_DFF2(.CK(recv_CK), .D(hrecv_G2), .Q(recv_G2), .SI(recv_G1), .SE(scan_enable));
SDFFNSR RECV_O_DFF0(.CK(recv_CK), .D(recv_G117), .Q(hrecv_G117), .SI(recv_G2), .SE(scan_enable));
SDFFNSR RECV_O_DFF1(.CK(recv_CK), .D(recv_G132), .Q(hrecv_G132), .SI(hrecv_G117), .SE(scan_enable));
SDFFNSR RECV_O_DFF2(.CK(recv_CK), .D(recv_G66), .Q(hrecv_G66), .SI(hrecv_G132), .SE(scan_enable));
SDFFNSR RECV_O_DFF3(.CK(recv_CK), .D(recv_G118), .Q(hrecv_G118), .SI(hrecv_G66), .SE(scan_enable));
SDFFNSR RECV_O_DFF4(.CK(recv_CK), .D(recv_G133), .Q(hrecv_G133), .SI(hrecv_G118), .SE(scan_enable));
SDFFNSR RECV_O_DFF5(.CK(recv_CK), .D(recv_G67), .Q(hrecv_G67), .SI(hrecv_G133), .SE(scan_enable));
// All orignal DFFs are extended into 2 copies
SDFFNSR SEND_DFF_0 (.CK(send_CK), .D(send_G29), .Q(send_G10), .SI(hrecv_G67), .SE(scan_enable));
SDFFNSR SEND_DFF_1 (.CK(send_CK), .D(send_G30), .Q(send_G11), .SI(send_G10), .SE(scan_enable));
SDFFNSR SEND_DFF_2 (.CK(send_CK), .D(send_G34), .Q(send_G12), .SI(send_G11), .SE(scan_enable));
SDFFNSR SEND_DFF_3 (.CK(send_CK), .D(send_G39), .Q(send_G13), .SI(send_G12), .SE(scan_enable));
SDFFNSR SEND_DFF_4 (.CK(send_CK), .D(send_G44), .Q(send_G14), .SI(send_G13), .SE(scan_enable));
SDFFNSR SEND_DFF_5 (.CK(send_CK), .D(send_G56), .Q(send_G15), .SI(send_G14), .SE(scan_enable));
SDFFNSR SEND_DFF_6 (.CK(send_CK), .D(send_G86), .Q(send_G16), .SI(send_G15), .SE(scan_enable));
SDFFNSR SEND_DFF_7 (.CK(send_CK), .D(send_G92), .Q(send_G17), .SI(send_G16), .SE(scan_enable));
SDFFNSR SEND_DFF_8 (.CK(send_CK), .D(send_G98), .Q(send_G18), .SI(send_G17), .SE(scan_enable));
SDFFNSR SEND_DFF_9 (.CK(send_CK), .D(send_G102), .Q(send_G19), .SI(send_G18), .SE(scan_enable));
SDFFNSR SEND_DFF_10 (.CK(send_CK), .D(send_G107), .Q(send_G20), .SI(send_G19), .SE(scan_enable));
SDFFNSR SEND_DFF_11 (.CK(send_CK), .D(send_G113), .Q(send_G21), .SI(send_G20), .SE(scan_enable));
SDFFNSR SEND_DFF_12 (.CK(send_CK), .D(send_G119), .Q(send_G22), .SI(send_G21), .SE(scan_enable));
SDFFNSR SEND_DFF_13 (.CK(send_CK), .D(send_G125), .Q(send_G23), .SI(send_G22), .SE(scan_enable));
SDFFNSR RECV_DFF_0 (.CK(recv_CK), .D(recv_G29), .Q(recv_G10), .SI(send_G23), .SE(scan_enable));
SDFFNSR RECV_DFF_1 (.CK(recv_CK), .D(recv_G30), .Q(recv_G11), .SI(recv_G10), .SE(scan_enable));
SDFFNSR RECV_DFF_2 (.CK(recv_CK), .D(recv_G34), .Q(recv_G12), .SI(recv_G11), .SE(scan_enable));
SDFFNSR RECV_DFF_3 (.CK(recv_CK), .D(recv_G39), .Q(recv_G13), .SI(recv_G12), .SE(scan_enable));
SDFFNSR RECV_DFF_4 (.CK(recv_CK), .D(recv_G44), .Q(recv_G14), .SI(recv_G13), .SE(scan_enable));
SDFFNSR RECV_DFF_5 (.CK(recv_CK), .D(recv_G56), .Q(recv_G15), .SI(recv_G14), .SE(scan_enable));
SDFFNSR RECV_DFF_6 (.CK(recv_CK), .D(recv_G86), .Q(recv_G16), .SI(recv_G15), .SE(scan_enable));
SDFFNSR RECV_DFF_7 (.CK(recv_CK), .D(recv_G92), .Q(recv_G17), .SI(recv_G16), .SE(scan_enable));
SDFFNSR RECV_DFF_8 (.CK(recv_CK), .D(recv_G98), .Q(recv_G18), .SI(recv_G17), .SE(scan_enable));
SDFFNSR RECV_DFF_9 (.CK(recv_CK), .D(recv_G102), .Q(recv_G19), .SI(recv_G18), .SE(scan_enable));
SDFFNSR RECV_DFF_10 (.CK(recv_CK), .D(recv_G107), .Q(recv_G20), .SI(recv_G19), .SE(scan_enable));
SDFFNSR RECV_DFF_11 (.CK(recv_CK), .D(recv_G113), .Q(recv_G21), .SI(recv_G20), .SE(scan_enable));
SDFFNSR RECV_DFF_12 (.CK(recv_CK), .D(recv_G119), .Q(recv_G22), .SI(recv_G21), .SE(scan_enable));
SDFFNSR RECV_DFF_13 (.CK(recv_CK), .D(recv_G125), .Q(recv_G23), .SI(recv_G22), .SE(scan_enable));
//END: All orignal DFFs are extended into 2 copies// scan chain ends here

buf1 BUF(scan_data_out, recv_G23);

not SEND_NOT_0(send_G28, send_G130);
not RECV_NOT_0(recv_G28, recv_G130);
not SEND_NOT_1(send_G38, send_G10);
not RECV_NOT_1(recv_G38, recv_G10);
not SEND_NOT_2(send_G40, send_G13);
not RECV_NOT_2(recv_G40, recv_G13);
not SEND_NOT_3(send_G45, send_G12);
not RECV_NOT_3(recv_G45, recv_G12);
not SEND_NOT_4(send_G46, send_G11);
not RECV_NOT_4(recv_G46, recv_G11);
not SEND_NOT_5(send_G50, send_G14);
not RECV_NOT_5(recv_G50, recv_G14);
not SEND_NOT_6(send_G51, send_G23);
not RECV_NOT_6(recv_G51, recv_G23);
not SEND_NOT_7(send_G54, send_G11);
not RECV_NOT_7(recv_G54, recv_G11);
not SEND_NOT_8(send_G55, send_G13);
not RECV_NOT_8(recv_G55, recv_G13);
not SEND_NOT_9(send_G59, send_G12);
not RECV_NOT_9(recv_G59, recv_G12);
not SEND_NOT_10(send_G60, send_G22);
not RECV_NOT_10(recv_G60, recv_G22);
not SEND_NOT_11(send_G64, send_G15);
not RECV_NOT_11(recv_G64, recv_G15);
not SEND_NOT_12(send_II155, send_G16);
not RECV_NOT_12(recv_II155, recv_G16);
not SEND_NOT_13(send_G66, send_II155);
not RECV_NOT_13(recv_G66, recv_II155);
not SEND_NOT_14(send_II158, send_G17);
not RECV_NOT_14(recv_II158, recv_G17);
not SEND_NOT_15(send_G67, send_II158);
not RECV_NOT_15(recv_G67, recv_II158);
not SEND_NOT_16(send_G76, send_G10);
not RECV_NOT_16(recv_G76, recv_G10);
not SEND_NOT_17(send_G82, send_G11);
not RECV_NOT_17(recv_G82, recv_G11);
not SEND_NOT_18(send_G87, send_G16);
not RECV_NOT_18(recv_G87, recv_G16);
not SEND_NOT_19(send_G91, send_G12);
not RECV_NOT_19(recv_G91, recv_G12);
not SEND_NOT_20(send_G93, send_G17);
not RECV_NOT_20(recv_G93, recv_G17);
not SEND_NOT_21(send_G96, send_G14);
not RECV_NOT_21(recv_G96, recv_G14);
not SEND_NOT_22(send_G99, send_G18);
not RECV_NOT_22(recv_G99, recv_G18);
not SEND_NOT_23(send_G103, send_G13);
not RECV_NOT_23(recv_G103, recv_G13);
not SEND_NOT_24(send_G108, send_G112);
not RECV_NOT_24(recv_G108, recv_G112);
not SEND_NOT_25(send_G114, send_G21);
not RECV_NOT_25(recv_G114, recv_G21);
not SEND_NOT_26(send_II210, send_G18);
not RECV_NOT_26(recv_II210, recv_G18);
not SEND_NOT_27(send_G117, send_II210);
not RECV_NOT_27(recv_G117, recv_II210);
not SEND_NOT_28(send_II213, send_G19);
not RECV_NOT_28(recv_II213, recv_G19);
not SEND_NOT_29(send_G118, send_II213);
not RECV_NOT_29(recv_G118, recv_II213);
not SEND_NOT_30(send_G120, send_G124);
not RECV_NOT_30(recv_G120, recv_G124);
not SEND_NOT_31(send_G121, send_G22);
not RECV_NOT_31(recv_G121, recv_G22);
not SEND_NOT_32(send_II221, send_G2);
not RECV_NOT_32(recv_II221, recv_G2);
not SEND_NOT_33(send_G124, send_II221);
not RECV_NOT_33(recv_G124, recv_II221);
not SEND_NOT_34(send_G126, send_G131);
not RECV_NOT_34(recv_G126, recv_G131);
not SEND_NOT_35(send_G127, send_G23);
not RECV_NOT_35(recv_G127, recv_G23);
not SEND_NOT_36(send_II229, send_G0);
not RECV_NOT_36(recv_II229, recv_G0);
not SEND_NOT_37(send_G130, send_II229);
not RECV_NOT_37(recv_G130, recv_II229);
not SEND_NOT_38(send_II232, send_G1);
not RECV_NOT_38(recv_II232, recv_G1);
not SEND_NOT_39(send_G131, send_II232);
not RECV_NOT_39(recv_G131, recv_II232);
not SEND_NOT_40(send_II235, send_G20);
not RECV_NOT_40(recv_II235, recv_G20);
not SEND_NOT_41(send_G132, send_II235);
not RECV_NOT_41(recv_G132, recv_II235);
not SEND_NOT_42(send_II238, send_G21);
not RECV_NOT_42(recv_II238, recv_G21);
not SEND_NOT_43(send_G133, send_II238);
not RECV_NOT_43(recv_G133, recv_II238);
and SEND_AND2_0(send_G26, send_G28, send_G50);
and RECV_AND2_0(recv_G26, recv_G28, recv_G50);
and SEND_AND2_1(send_G27, send_G51, send_G28);
and RECV_AND2_1(recv_G27, recv_G51, recv_G28);
and SEND_AND3_0(send_G31, send_G10, send_G45, send_G13);
and RECV_AND3_0(recv_G31, recv_G10, recv_G45, recv_G13);
and SEND_AND2_2(send_G32, send_G10, send_G11);
and RECV_AND2_2(recv_G32, recv_G10, recv_G11);
and SEND_AND2_3(send_G33, send_G38, send_G46);
and RECV_AND2_3(recv_G33, recv_G38, recv_G46);
and SEND_AND3_1(send_G35, send_G10, send_G11, send_G12);
and RECV_AND3_1(recv_G35, recv_G10, recv_G11, recv_G12);
and SEND_AND2_4(send_G36, send_G38, send_G45);
and RECV_AND2_4(recv_G36, recv_G38, recv_G45);
and SEND_AND2_5(send_G37, send_G46, send_G45);
and RECV_AND2_5(recv_G37, recv_G46, recv_G45);
and SEND_AND2_6(send_G42, send_G40, send_G41);
and RECV_AND2_6(recv_G42, recv_G40, recv_G41);
and SEND_AND4_0(send_G48, send_G45, send_G46, send_G10, send_G47);
and RECV_AND4_0(recv_G48, recv_G45, recv_G46, recv_G10, recv_G47);
and SEND_AND3_2(send_G49, send_G50, send_G51, send_G52);
and RECV_AND3_2(recv_G49, recv_G50, recv_G51, recv_G52);
and SEND_AND4_1(send_G57, send_G59, send_G11, send_G60, send_G61);
and RECV_AND4_1(recv_G57, recv_G59, recv_G11, recv_G60, recv_G61);
and SEND_AND2_7(send_G58, send_G64, send_G65);
and RECV_AND2_7(recv_G58, recv_G64, recv_G65);
and SEND_AND4_2(send_G62, send_G59, send_G11, send_G60, send_G61);
and RECV_AND4_2(recv_G62, recv_G59, recv_G11, recv_G60, recv_G61);
and SEND_AND2_8(send_G63, send_G64, send_G65);
and RECV_AND2_8(recv_G63, recv_G64, recv_G65);
and SEND_AND3_3(send_G74, send_G12, send_G14, send_G19);
and RECV_AND3_3(recv_G74, recv_G12, recv_G14, recv_G19);
and SEND_AND3_4(send_G75, send_G82, send_G91, send_G14);
and RECV_AND3_4(recv_G75, recv_G82, recv_G91, recv_G14);
and SEND_AND2_9(send_G88, send_G14, send_G87);
and RECV_AND2_9(recv_G88, recv_G14, recv_G87);
and SEND_AND2_10(send_G89, send_G103, send_G96);
and RECV_AND2_10(recv_G89, recv_G103, recv_G96);
and SEND_AND2_11(send_G90, send_G91, send_G103);
and RECV_AND2_11(recv_G90, recv_G91, recv_G103);
and SEND_AND2_12(send_G94, send_G93, send_G13);
and RECV_AND2_12(recv_G94, recv_G93, recv_G13);
and SEND_AND2_13(send_G95, send_G96, send_G13);
and RECV_AND2_13(recv_G95, recv_G96, recv_G13);
and SEND_AND3_5(send_G100, send_G99, send_G14, send_G12);
and RECV_AND3_5(recv_G100, recv_G99, recv_G14, recv_G12);
and SEND_AND3_6(send_G105, send_G103, send_G108, send_G104);
and RECV_AND3_6(recv_G105, recv_G103, recv_G108, recv_G104);
and SEND_AND2_14(send_G110, send_G108, send_G109);
and RECV_AND2_14(recv_G110, recv_G108, recv_G109);
and SEND_AND2_15(send_G111, send_G10, send_G112);
and RECV_AND2_15(recv_G111, recv_G10, recv_G112);
and SEND_AND2_16(send_G115, send_G114, send_G14);
and RECV_AND2_16(recv_G115, recv_G114, recv_G14);
and SEND_AND2_17(send_G122, send_G120, send_G121);
and RECV_AND2_17(recv_G122, recv_G120, recv_G121);
and SEND_AND2_18(send_G123, send_G124, send_G22);
and RECV_AND2_18(recv_G123, recv_G124, recv_G22);
and SEND_AND2_19(send_G128, send_G126, send_G127);
and RECV_AND2_19(recv_G128, recv_G126, recv_G127);
and SEND_AND2_20(send_G129, send_G131, send_G23);
and RECV_AND2_20(recv_G129, recv_G131, recv_G23);
or SEND_OR4_0(send_G24, send_G38, send_G46, send_G45, send_G40);
or RECV_OR4_0(recv_G24, recv_G38, recv_G46, recv_G45, recv_G40);
or SEND_OR3_0(send_G25, send_G38, send_G11, send_G12);
or RECV_OR3_0(recv_G25, recv_G38, recv_G11, recv_G12);
or SEND_OR4_1(send_G68, send_G11, send_G12, send_G13, send_G96);
or RECV_OR4_1(recv_G68, recv_G11, recv_G12, recv_G13, recv_G96);
or SEND_OR2_0(send_G69, send_G103, send_G18);
or RECV_OR2_0(recv_G69, recv_G103, recv_G18);
or SEND_OR2_1(send_G70, send_G103, send_G14);
or RECV_OR2_1(recv_G70, recv_G103, recv_G14);
or SEND_OR3_1(send_G71, send_G82, send_G12, send_G13);
or RECV_OR3_1(recv_G71, recv_G82, recv_G12, recv_G13);
or SEND_OR2_2(send_G72, send_G91, send_G20);
or RECV_OR2_2(recv_G72, recv_G91, recv_G20);
or SEND_OR2_3(send_G73, send_G103, send_G20);
or RECV_OR2_3(recv_G73, recv_G103, recv_G20);
or SEND_OR4_2(send_G77, send_G112, send_G103, send_G96, send_G19);
or RECV_OR4_2(recv_G77, recv_G112, recv_G103, recv_G96, recv_G19);
or SEND_OR2_4(send_G78, send_G108, send_G76);
or RECV_OR2_4(recv_G78, recv_G108, recv_G76);
or SEND_OR2_5(send_G79, send_G103, send_G14);
or RECV_OR2_5(recv_G79, recv_G103, recv_G14);
or SEND_OR2_6(send_G80, send_G11, send_G14);
or RECV_OR2_6(recv_G80, recv_G11, recv_G14);
or SEND_OR2_7(send_G81, send_G12, send_G13);
or RECV_OR2_7(recv_G81, recv_G12, recv_G13);
or SEND_OR4_3(send_G83, send_G11, send_G12, send_G13, send_G96);
or RECV_OR4_3(recv_G83, recv_G11, recv_G12, recv_G13, recv_G96);
or SEND_OR3_2(send_G84, send_G82, send_G91, send_G14);
or RECV_OR3_2(recv_G84, recv_G82, recv_G91, recv_G14);
or SEND_OR3_3(send_G85, send_G91, send_G96, send_G17);
or RECV_OR3_3(recv_G85, recv_G91, recv_G96, recv_G17);
nand SEND_NAND3_0(send_G41, send_G12, send_G11, send_G10);
nand RECV_NAND3_0(recv_G41, recv_G12, recv_G11, recv_G10);
nand SEND_NAND3_1(send_G43, send_G24, send_G25, send_G28);
nand RECV_NAND3_1(recv_G43, recv_G24, recv_G25, recv_G28);
nand SEND_NAND4_0(send_G52, send_G13, send_G45, send_G46, send_G10);
nand RECV_NAND4_0(recv_G52, recv_G13, recv_G45, recv_G46, recv_G10);
nand SEND_NAND4_1(send_G65, send_G59, send_G54, send_G22, send_G61);
nand RECV_NAND4_1(recv_G65, recv_G59, recv_G54, recv_G22, recv_G61);
nand SEND_NAND4_2(send_G97, send_G83, send_G84, send_G85, send_G108);
nand RECV_NAND4_2(recv_G97, recv_G83, recv_G84, recv_G85, recv_G108);
nand SEND_NAND4_3(send_G101, send_G68, send_G69, send_G70, send_G108);
nand RECV_NAND4_3(recv_G101, recv_G68, recv_G69, recv_G70, recv_G108);
nand SEND_NAND2_0(send_G106, send_G77, send_G78);
nand RECV_NAND2_0(recv_G106, recv_G77, recv_G78);
nand SEND_NAND4_4(send_G109, send_G71, send_G72, send_G73, send_G14);
nand RECV_NAND4_4(recv_G109, recv_G71, recv_G72, recv_G73, recv_G14);
nand SEND_NAND4_5(send_G116, send_G79, send_G80, send_G81, send_G108);
nand RECV_NAND4_5(recv_G116, recv_G79, recv_G80, recv_G81, recv_G108);
nor SEND_NOR2_0(send_G29, send_G10, send_G130);
nor RECV_NOR2_0(recv_G29, recv_G10, recv_G130);
nor SEND_NOR4_0(send_G30, send_G31, send_G32, send_G33, send_G130);
nor RECV_NOR4_0(recv_G30, recv_G31, recv_G32, recv_G33, recv_G130);
nor SEND_NOR4_1(send_G34, send_G35, send_G36, send_G37, send_G130);
nor RECV_NOR4_1(recv_G34, recv_G35, recv_G36, recv_G37, recv_G130);
nor SEND_NOR2_1(send_G39, send_G42, send_G43);
nor RECV_NOR2_1(recv_G39, recv_G42, recv_G43);
nor SEND_NOR3_0(send_G44, send_G48, send_G49, send_G53);
nor RECV_NOR3_0(recv_G44, recv_G48, recv_G49, recv_G53);
nor SEND_NOR2_2(send_G47, send_G50, send_G40);
nor RECV_NOR2_2(recv_G47, recv_G50, recv_G40);
nor SEND_NOR2_3(send_G53, send_G26, send_G27);
nor RECV_NOR2_3(recv_G53, recv_G26, recv_G27);
nor SEND_NOR3_1(send_G56, send_G57, send_G58, send_G130);
nor RECV_NOR3_1(recv_G56, recv_G57, recv_G58, recv_G130);
nor SEND_NOR2_4(send_G61, send_G14, send_G55);
nor RECV_NOR2_4(recv_G61, recv_G14, recv_G55);
nor SEND_NOR4_2(send_G86, send_G88, send_G89, send_G90, send_G112);
nor RECV_NOR4_2(recv_G86, recv_G88, recv_G89, recv_G90, recv_G112);
nor SEND_NOR3_2(send_G92, send_G94, send_G95, send_G97);
nor RECV_NOR3_2(recv_G92, recv_G94, recv_G95, recv_G97);
nor SEND_NOR2_5(send_G98, send_G100, send_G101);
nor RECV_NOR2_5(recv_G98, recv_G100, recv_G101);
nor SEND_NOR2_6(send_G102, send_G105, send_G106);
nor RECV_NOR2_6(recv_G102, recv_G105, recv_G106);
nor SEND_NOR2_7(send_G104, send_G74, send_G75);
nor RECV_NOR2_7(recv_G104, recv_G74, recv_G75);
nor SEND_NOR2_8(send_G107, send_G110, send_G111);
nor RECV_NOR2_8(recv_G107, recv_G110, recv_G111);
nor SEND_NOR2_9(send_G112, send_G62, send_G63);
nor RECV_NOR2_9(recv_G112, recv_G62, recv_G63);
nor SEND_NOR2_10(send_G113, send_G115, send_G116);
nor RECV_NOR2_10(recv_G113, recv_G115, recv_G116);
nor SEND_NOR3_3(send_G119, send_G122, send_G123, send_G130);
nor RECV_NOR3_3(recv_G119, recv_G122, recv_G123, recv_G130);
nor SEND_NOR3_4(send_G125, send_G128, send_G129, send_G130);
nor RECV_NOR3_4(recv_G125, recv_G128, recv_G129, recv_G130);
endmodule

module buf1 (out, in);
    output out;
    input in;
    buf (out, in);
endmodule
    

//# 46 DFFs