
module buf1 (out, in);
    output out;
    input in;
    buf (out, in);
endmodule
    module bit_clk_pad_i_domain (scan_enable, scan_data_in, scan_data_out, bit_clk_pad_i, out_slt3, out_slt_67, out_slt_146, out_slt_102, out_slt_175, out_slt_168, crac_out_867, crac_out_876, crac_out_866, out_slt_145, crac_out_848, out_slt_162, out_slt_129, crac_out_858, out_slt_20, out_slt_19, out_slt_18, out_slt_80, out_slt_164, crac_out_846, out_slt_158, out_slt_77, out_slt_143, out_slt_166, crac_out_850, out_slt_73, out_slt_81, crac_out_856, out_slt_66, out_slt_173, out_slt_78, out_slt6, out_slt_136, out_slt_123, out_slt_161, out_slt_101, out_slt_128, out_slt_157, crac_out_859, out_slt_178, out_slt_138, out_slt_121, out_slt_83, out_slt_169, out_slt_156, crac_out_857, out_slt_110, crac_out_860, out_slt_74, out_slt_113, out_slt_170, out_slt_122, crac_out_849, out_slt_72, out_slt_115, out_slt_65, out_slt_159, out_slt_108, out_slt_105, out_slt4, out_slt_96, u1_sdata_in_r, out_slt_167, out_slt_127, out_slt_176, out_slt_140, crac_out_847, out_slt_165, out_slt_117, out_slt_95, out_slt_93, crac_out, out_slt_120, out_slt_76, out_slt_126, out_slt_131, out_slt_139, crac_out_851, out_slt_142, crac_out_854, out_slt_135, out_slt_151, out_slt_137, out_slt_132, out_slt_22, out_slt_23, out_slt_24, out_slt_25, out_slt_125, crac_out_852, out_slt_171, out_slt_153, out_slt_144, crac_out_864, crac_out_865, crac_out_862, crac_out_863, crac_out_861, out_slt7, out_slt_152, out_slt_104, out_slt_91, out_slt_82, out_slt_130, suspended_o, out_slt_119, out_slt_174, out_slt_155, out_slt_154, out_slt_147, out_slt_87, crac_out_855, out_slt_98, out_slt_172, out_slt8, out_slt_133, out_slt_75, out_slt_92, out_slt_114, out_slt_106, out_slt_124, out_slt_100, out_slt_17, out_slt_160, out_slt_85, out_slt_79, out_slt_116, out_slt_71, out_slt_89, out_slt_84, out_slt_148, out_slt_70, out_slt_111, out_slt_99, out_slt_86, out_slt_103, out_slt_118, out_slt_107, out_slt_150, out_slt_97, crac_out_853, out_slt_112, out_slt_94, out_slt_88, out_slt_69, out_slt9, out_slt_177, out_slt_134, out_slt_141, out_slt_163, out_slt_90, out_slt_149, out_slt_68, out_slt_109, in_valid_9, u2_sync_beat, in_valid, valid, sdata_pad_o);

input scan_enable, scan_data_in, bit_clk_pad_i, out_slt3, out_slt_67, out_slt_146, out_slt_102, out_slt_175, out_slt_168, crac_out_867, crac_out_876, crac_out_866, out_slt_145, crac_out_848, out_slt_162, out_slt_129, crac_out_858, out_slt_20, out_slt_19, out_slt_18, out_slt_80, out_slt_164, crac_out_846, out_slt_158, out_slt_77, out_slt_143, out_slt_166, crac_out_850, out_slt_73, out_slt_81, crac_out_856, out_slt_66, out_slt_173, out_slt_78, out_slt6, out_slt_136, out_slt_123, out_slt_161, out_slt_101, out_slt_128, out_slt_157, crac_out_859, out_slt_178, out_slt_138, out_slt_121, out_slt_83, out_slt_169, out_slt_156, crac_out_857, out_slt_110, crac_out_860, out_slt_74, out_slt_113, out_slt_170, out_slt_122, crac_out_849, out_slt_72, out_slt_115, out_slt_65, out_slt_159, out_slt_108, out_slt_105, out_slt4, out_slt_96, u1_sdata_in_r, out_slt_167, out_slt_127, out_slt_176, out_slt_140, crac_out_847, out_slt_165, out_slt_117, out_slt_95, out_slt_93, crac_out, out_slt_120, out_slt_76, out_slt_126, out_slt_131, out_slt_139, crac_out_851, out_slt_142, crac_out_854, out_slt_135, out_slt_151, out_slt_137, out_slt_132, out_slt_22, out_slt_23, out_slt_24, out_slt_25, out_slt_125, crac_out_852, out_slt_171, out_slt_153, out_slt_144, crac_out_864, crac_out_865, crac_out_862, crac_out_863, crac_out_861, out_slt7, out_slt_152, out_slt_104, out_slt_91, out_slt_82, out_slt_130, suspended_o, out_slt_119, out_slt_174, out_slt_155, out_slt_154, out_slt_147, out_slt_87, crac_out_855, out_slt_98, out_slt_172, out_slt8, out_slt_133, out_slt_75, out_slt_92, out_slt_114, out_slt_106, out_slt_124, out_slt_100, out_slt_17, out_slt_160, out_slt_85, out_slt_79, out_slt_116, out_slt_71, out_slt_89, out_slt_84, out_slt_148, out_slt_70, out_slt_111, out_slt_99, out_slt_86, out_slt_103, out_slt_118, out_slt_107, out_slt_150, out_slt_97, crac_out_853, out_slt_112, out_slt_94, out_slt_88, out_slt_69, out_slt9, out_slt_177, out_slt_134, out_slt_141, out_slt_163, out_slt_90, out_slt_149, out_slt_68, out_slt_109;
output scan_data_out, in_valid_9, u2_sync_beat, in_valid, valid, sdata_pad_o;
wire n_11214;
wire n_208;
wire u0_slt9_r_182;
wire n_11395;
wire n_11213;
wire n_297;
wire u0_slt9_r_181;
wire n_11319;
wire n_11312;
wire n_10790;
wire u0_slt4_r_73;
wire n_6710;
wire n_11211;
wire n_203;
wire u0_slt9_r_179;
wire n_11389;
wire n_11314;
wire n_373;
wire u0_slt4_r_75;
wire n_11313;
wire n_10788;
wire u0_slt4_r_74;
wire n_11317;
wire n_370;
wire u0_slt4_r_77;
wire n_11315;
wire n_380;
wire u0_slt4_r_76;
wire n_7042;
wire in_slt_739;
wire n_9958;
wire n_866;
wire n_5821;
wire n_698;
wire u2_cnt_b3_b;
wire u0_slt6_r_117;
wire n_11272;
wire u0_slt1_r_34;
wire n_11417;
wire in_slt_426;
wire n_9354;
wire in_slt_402;
wire n_7509;
wire n_11212;
wire n_263;
wire u0_slt9_r_180;
wire n_11210;
wire n_152;
wire u0_slt9_r_178;
wire in_slt_425;
wire n_8255;
wire u1_sr_120;
wire u1_sr_119;
wire n_1928;
wire n_688;
wire n_1824;
wire n_5430;
wire n_2572;
wire u2_cnt_b6_b;
wire n_1212;
wire in_slt_409;
wire n_10803;
wire in_slt_444;
wire n_7154;
wire n_4840;
wire in_slt_455;
wire n_11114;
wire n_251;
wire u0_slt9_r_177;
wire n_11207;
wire u0_slt7_r_141;
wire n_11253;
wire u0_slt5_r_103;
wire n_11301;
wire u0_slt9_r_185;
wire n_11216;
wire n_11243;
wire n_10990;
wire u0_slt7_r_130;
wire n_11246;
wire n_201;
wire u0_slt7_r_133;
wire n_11247;
wire n_217;
wire u0_slt7_r_134;
wire n_11244;
wire n_10988;
wire u0_slt7_r_131;
wire n_11245;
wire n_335;
wire u0_slt7_r_132;
wire u0_slt1_r_26;
wire n_11406;
wire u0_slt7_r_148;
wire n_11262;
wire in_slt_450;
wire n_9618;
wire u1_sr_126;
wire u1_sr_125;
wire n_10976;
wire n_352;
wire n_361;
wire in_slt_748;
wire n_7507;
wire n_5741;
wire n_4826;
wire n_6057;
wire u1_sr_135;
wire u1_sr_134;
wire u0_slt5_r_93;
wire n_11291;
wire n_4107;
wire n_1823;
wire n_1469;
wire n_7043;
wire n_1087;
wire in_slt_433;
wire n_11115;
wire u0_slt2_r_43;
wire n_11376;
wire u0_slt4_r_78;
wire u0_slt2_r_53;
wire n_11390;
wire u0_slt2_r_50;
wire n_11385;
wire u0_slt3_r_63;
wire n_11351;
wire n_183;
wire u1_sr_118;
wire u0_slt6_r_120;
wire n_11276;
wire n_11235;
wire n_228;
wire u0_slt8_r_161;
wire n_11234;
wire n_76;
wire u0_slt8_r_160;
wire n_11237;
wire n_79;
wire u0_slt8_r_163;
wire n_11236;
wire n_237;
wire u0_slt8_r_162;
wire n_11233;
wire n_212;
wire u0_slt8_r_159;
wire u0_slt9_r_168;
wire n_8211;
wire u0_slt6_r_128;
wire n_11287;
wire u1_sr_128;
wire out_le;
wire n_11416;
wire u0_slt1_r_32;
wire u0_slt1_r_33;
wire n_11418;
wire n_11419;
wire u0_slt0_r;
wire n_11414;
wire u0_slt1_r_31;
wire n_11258;
wire n_163;
wire u0_slt7_r_145;
wire n_299;
wire u0_slt7_r_147;
wire u0_slt4_r_79;
wire n_11318;
wire u0_slt9_r_176;
wire n_11206;
wire in_slt_749;
wire n_8258;
wire u0_slt8_r_154;
wire n_11225;
wire u0_slt1_r_22;
wire n_11400;
wire u0_slt3_r_56;
wire n_11341;
wire u0_slt1_r;
wire n_11391;
wire n_280;
wire n_7038;
wire n_6734;
wire n_71;
wire in_slt_404;
wire n_9355;
wire u0_slt1_r_23;
wire n_11401;
wire u0_slt5_r_102;
wire n_11303;
wire u0_slt5_r_104;
wire n_11302;
wire n_11305;
wire u0_slt5_r_106;
wire n_11304;
wire u0_slt5_r_105;
wire in_slt_397;
wire n_6732;
wire n_2597;
wire n_9619;
wire in_slt_428;
wire out_le_183;
wire n_9625;
wire in_slt_406;
wire out_le_182;
wire n_9952;
wire n_265;
wire n_179;
wire n_6721;
wire in_slt_443;
wire out_le_184;
wire n_6722;
wire in_slt_442;
wire n_6728;
wire u1_sr;
wire in_slt4;
wire n_7358;
wire u1_sr_121;
wire in_slt_401;
wire n_6726;
wire in_slt_420;
wire n_6727;
wire u1_sr_117;
wire in_slt_419;
wire n_7155;
wire in_slt_422;
wire n_6723;
wire in_slt_441;
wire in_slt_838;
wire n_9957;
wire n_1825;
wire n_1822;
wire n_684;
wire n_11431;
wire u0_slt0_r_9;
wire n_11430;
wire u0_slt0_r_8;
wire n_11429;
wire u0_slt0_r_7;
wire n_11428;
wire u0_slt0_r_6;
wire n_5611;
wire n_3965;
wire n_3995;
wire n_4079;
wire u0_slt4_r_84;
wire n_11326;
wire n_11427;
wire n_281;
wire n_359;
wire n_11205;
wire n_160;
wire u0_slt9_r_174;
wire u0_slt9_r_175;
wire n_5889;
wire n_11307;
wire u0_slt5_r_108;
wire n_11308;
wire u0_slt5_r_109;
wire n_5593;
wire in_slt_845;
wire n_11202;
wire n_6999;
wire u0_slt0_r_5;
wire n_11424;
wire u0_slt6_r_112;
wire n_11266;
wire n_11292;
wire n_11293;
wire u0_slt5_r_94;
wire n_11294;
wire u0_slt5_r_95;
wire n_11295;
wire u0_slt5_r_96;
wire u0_slt5_r_92;
wire n_227;
wire n_86;
wire n_5441;
wire n_3996;
wire n_4832;
wire n_456;
wire n_701;
wire u2_cnt_b5_b;
wire n_4825;
wire n_4095;
wire n_11387;
wire n_11392;
wire n_11388;
wire n_177;
wire u0_slt2_r_51;
wire n_170;
wire u0_slt2_r_52;
wire n_11300;
wire u0_slt9_r_183;
wire n_195;
wire u1_sr_131;
wire u1_sr_130;
wire n_2632;
wire n_2631;
wire n_11284;
wire n_113;
wire u0_slt6_r_125;
wire n_11283;
wire n_101;
wire u0_slt6_r_124;
wire n_11166;
wire u1_sr_132;
wire in_slt_456;
wire n_11281;
wire n_261;
wire u0_slt6_r_123;
wire n_11280;
wire n_300;
wire u0_slt6_r_122;
wire n_11279;
wire n_84;
wire u0_slt6_r_121;
wire in_slt_430;
wire n_9955;
wire n_1785;
wire n_1784;
wire n_1782;
wire n_2592;
wire n_3964;
wire n_2596;
wire n_11200;
wire in_slt_437;
wire u0_slt2_r_38;
wire n_11370;
wire u0_slt4_r_81;
wire n_11321;
wire n_5635;
wire n_4103;
wire u0_slt7_r_140;
wire n_11252;
wire in_slt_753;
wire n_9764;
wire u0_slt2_r_47;
wire n_11381;
wire u0_slt1_r_25;
wire n_11404;
wire n_11203;
wire n_372;
wire u0_slt9_r_172;
wire in_slt_750;
wire n_9357;
wire n_11403;
wire u0_slt1_r_24;
wire u0_slt1_r_21;
wire u0_slt2_r_35;
wire n_11365;
wire n_1486;
wire u0_slt8_r_149;
wire n_11219;
wire n_1100;
wire n_10981;
wire n_191;
wire u0_slt3_r_57;
wire n_11342;
wire u1_sr_123;
wire out_le_180;
wire u0_slt3_r_70;
wire n_11360;
wire n_10785;
wire u0_slt6_r_111;
wire n_11269;
wire n_262;
wire u0_slt6_r_114;
wire n_11270;
wire n_234;
wire u0_slt6_r_115;
wire n_11267;
wire n_10783;
wire n_11268;
wire n_304;
wire u0_slt6_r_113;
wire u0_slt6_r;
wire n_11263;
wire n_311;
wire u0_slt9_r_169;
wire n_9603;
wire n_7508;
wire u1_sr_122;
wire in_slt_446;
wire in_slt_436;
wire n_11196;
wire u0_slt8_r_164;
wire n_2571;
wire u0_slt1_r_16;
wire in_slt_405;
wire n_9529;
wire u0_slt4_r_89;
wire n_11332;
wire u0_slt7_r_137;
wire n_11249;
wire u0_slt4_r_82;
wire n_11323;
wire u0_slt4_r_90;
wire n_11333;
wire n_341;
wire u2_cnt_b2_b;
wire n_109;
wire in_slt_398;
wire n_6730;
wire n_138;
wire n_10978;
wire n_2602;
wire n_2603;
wire in_slt_839;
wire n_10804;
wire n_10957;
wire in_slt_454;
wire n_10964;
wire in_slt_840;
wire out_le_181;
wire n_10958;
wire in_slt_432;
wire n_10961;
wire in_slt_410;
wire u1_sr_124;
wire n_11373;
wire u0_slt2_r_40;
wire u0_slt5_r;
wire n_11289;
wire n_11378;
wire n_357;
wire u0_slt2_r_44;
wire n_11377;
wire n_149;
wire u0_slt2_r_42;
wire n_11375;
wire n_130;
wire u0_slt2_r_41;
wire n_11361;
wire n_16;
wire n_6066;
wire u0_slt5_r_100;
wire n_11298;
wire n_7510;
wire in_slt_832;
wire n_267;
wire n_4096;
wire n_223;
wire n_134;
wire n_394;
wire u0_slt4_r_80;
wire n_11320;
wire n_391;
wire n_11324;
wire n_321;
wire n_320;
wire n_351;
wire in_slt_411;
wire n_11116;
wire n_9602;
wire n_295;
wire n_363;
wire n_240;
wire in_slt_457;
wire n_11184;
wire u0_slt5_r_110;
wire n_383;
wire u0_slt0_r_14;
wire n_11436;
wire u0_slt7_r_143;
wire n_11255;
wire u0_slt5_r_101;
wire n_11299;
wire n_1253;
wire n_1227;
wire u2_cnt_b4_b;
wire n_11209;
wire n_9530;
wire in_slt_835;
wire n_9531;
wire in_slt_736;
wire n_9528;
wire in_slt_427;
wire n_3984;
wire n_2593;
wire in_slt_452;
wire n_9954;
wire u1_sr_127;
wire n_102;
wire n_329;
wire n_11311;
wire n_711;
wire in_slt_431;
wire n_10802;
wire n_396;
wire u0_slt4_r_88;
wire n_11334;
wire n_11336;
wire u0_slt4_r_91;
wire n_11338;
wire n_220;
wire u0_slt3_r;
wire n_308;
wire n_4833;
wire n_5432;
wire n_4000;
wire n_4831;
wire n_1114;
wire n_2604;
wire n_2378;
wire n_338;
wire u0_slt3_r_65;
wire n_11353;
wire n_266;
wire u0_slt3_r_72;
wire n_11363;
wire u1_sr_129;
wire u0_slt8_r_157;
wire n_11230;
wire n_1520;
wire u0_slt8_r;
wire n_11218;
wire n_11204;
wire n_1774;
wire n_1519;
wire n_1773;
wire u0_slt3_r_58;
wire n_11344;
wire u0_slt1_r_20;
wire n_11397;
wire n_7003;
wire n_389;
wire n_287;
wire n_302;
wire in_slt_831;
wire n_7360;
wire n_11347;
wire n_230;
wire u0_slt3_r_59;
wire n_11352;
wire n_398;
wire u0_slt3_r_62;
wire n_11349;
wire u0_slt3_r_61;
wire n_11348;
wire n_82;
wire u0_slt3_r_60;
wire n_22;
wire in_slt_399;
wire n_6729;
wire in_slt_844;
wire n_11198;
wire u0_slt7_r_135;
wire u0_slt7_r_138;
wire n_11250;
wire u0_slt6_r_119;
wire n_11274;
wire in_slt_423;
wire n_7362;
wire u0_slt4_r_83;
wire n_328;
wire n_11364;
wire u0_slt2_r;
wire u0_slt3_r_71;
wire u0_slt3_r_69;
wire n_11242;
wire n_9628;
wire in_slt_836;
wire n_9630;
wire in_slt_752;
wire in_slt_414;
wire n_11197;
wire in_slt_449;
wire n_9527;
wire n_397;
wire n_330;
wire n_11290;
wire u0_slt0_r_11;
wire n_11433;
wire n_11306;
wire n_11010;
wire n_322;
wire u0_slt9_r_170;
wire n_11117;
wire in_slt_841;
wire n_11118;
wire in_slt_742;
wire n_150;
wire u0_slt7_r_142;
wire n_11254;
wire in_slt_747;
wire n_7359;
wire n_306;
wire n_11413;
wire u0_slt2_r_49;
wire n_11384;
wire u0_slt7_r_136;
wire n_375;
wire n_11251;
wire n_387;
wire n_229;
wire u0_slt7_r_139;
wire n_11248;
wire u0_slt4_r;
wire n_11310;
wire u0_slt6_r_127;
wire n_11286;
wire n_1213;
wire n_4076;
wire n_332;
wire u0_slt8_r_151;
wire n_11221;
wire n_11346;
wire u0_slt3_r_64;
wire u0_slt8_r_167;
wire n_11240;
wire in_slt_400;
wire n_7156;
wire n_392;
wire n_117;
wire u0_slt9_r;
wire n_7231;
wire n_157;
wire n_11399;
wire n_9763;
wire in_slt_837;
wire n_9762;
wire in_slt_407;
wire n_9761;
wire in_slt_429;
wire n_9765;
wire in_slt_738;
wire n_9760;
wire in_slt_451;
wire u0_slt4_r_87;
wire n_11329;
wire n_11217;
wire n_19;
wire u0_slt9_r_184;
wire n_57;
wire n_273;
wire u0_slt9_r_186;
wire n_11215;
wire n_1829;
wire n_6058;
wire n_6731;
wire in_slt3;
wire u0_slt6_r_118;
wire n_11273;
wire u0_slt5_r_97;
wire n_11368;
wire u0_slt2_r_36;
wire in_slt_421;
wire n_6725;
wire n_399;
wire n_9953;
wire n_9956;
wire in_slt_408;
wire in_slt6;
wire n_6724;
wire u0_slt5_r_107;
wire u0_slt9_r_173;
wire n_333;
wire in_slt_448;
wire n_9353;
wire in_slt_413;
wire n_11186;
wire n_674;
wire n_1355;
wire in_slt_459;
wire n_11199;
wire u0_slt0_r_12;
wire n_11434;
wire n_11257;
wire u0_slt2_r_45;
wire n_2629;
wire n_11366;
wire n_11423;
wire u0_slt0_r_3;
wire n_11238;
wire u0_slt7_r;
wire n_11241;
wire n_184;
wire u0_slt8_r_166;
wire n_11239;
wire u0_slt8_r_165;
wire u0_slt3_r_67;
wire n_11355;
wire u0_slt2_r_46;
wire n_11379;
wire n_11188;
wire n_11296;
wire n_11297;
wire u0_slt5_r_98;
wire u0_slt5_r_99;
wire n_10983;
wire u0_slt8_r_150;
wire n_11220;
wire n_11232;
wire n_112;
wire u0_slt1_r_18;
wire n_11394;
wire n_186;
wire n_181;
wire n_7144;
wire in_slt_830;
wire n_7361;
wire in_slt_445;
wire in_slt_833;
wire n_8257;
wire n_1552;
wire n_11231;
wire n_167;
wire u0_slt8_r_158;
wire n_11228;
wire n_376;
wire u0_slt8_r_155;
wire n_384;
wire u0_slt8_r_156;
wire n_11227;
wire n_362;
wire n_11421;
wire u0_slt0_r_2;
wire n_11425;
wire u0_slt0_r_4;
wire in_slt_834;
wire n_9356;
wire n_11420;
wire u0_slt0_r_1;
wire n_2377;
wire n_114;
wire u0_slt6_r_126;
wire u0_slt6_r_129;
wire n_11288;
wire n_1138;
wire n_11330;
wire n_254;
wire n_5820;
wire u0_slt6_r_116;
wire u0_slt0_r_10;
wire n_11435;
wire u0_slt0_r_13;
wire n_11437;
wire n_7013;
wire n_11438;
wire n_11426;
wire in_slt_447;
wire n_8254;
wire n_264;
wire n_166;
wire n_702;
wire n_11260;
wire n_11393;
wire in_slt_434;
wire n_11167;
wire u0_slt1_r_19;
wire n_11396;
wire u0_slt1_r_17;
wire u0_slt1_r_30;
wire n_11411;
wire u0_slt7_r_144;
wire n_11256;
wire n_11169;
wire in_slt_842;
wire n_11168;
wire in_slt_412;
wire u0_slt7_r_146;
wire n_11264;
wire n_21;
wire u0_slt2_r_39;
wire n_11371;
wire n_120;
wire n_11278;
wire n_182;
wire n_5448;
wire u0_slt8_r_153;
wire n_11224;
wire n_11201;
wire in_slt_415;
wire n_687;
wire u0_slt1_r_29;
wire n_11409;
wire u0_slt1_r_27;
wire n_11410;
wire u0_slt1_r_28;
wire n_11408;
wire u0_slt3_r_66;
wire n_11354;
wire n_11187;
wire u1_sr_133;
wire in_slt_843;
wire n_11185;
wire in_slt_435;
wire u0_slt4_r_85;
wire n_11327;
wire n_7511;
wire in_slt_424;
wire u0_slt9_r_171;
wire n_11195;
wire in_slt_458;
wire n_6052;
wire n_11328;
wire n_103;
wire n_243;
wire u0_slt4_r_86;
wire n_248;
wire n_56;
wire n_1372;
wire n_11383;
wire u0_slt2_r_48;
wire n_231;
wire n_401;
wire n_211;
wire n_200;
wire n_348;
wire u0_slt3_r_55;
wire n_11339;
wire u0_slt3_r_54;
wire n_11358;
wire n_7017;
wire n_11356;
wire n_282;
wire u0_slt3_r_68;
wire n_5822;
wire u0_slt8_r_152;
wire n_11223;
wire n_440;
wire n_679;
wire u0_slt2_r_37;
wire n_11372;
wire n_290;
wire n_1301;
wire n_4077;
wire in_slt_453;
wire n_10800;
wire n_1374;
wire n_8256;
wire in_slt_403;
wire n_259;
// scan chain begins here
SDFFNSRN u0_slt0_r_reg_b15_b (.CK(bit_clk_pad_i), .D(n_11438), .Q(sdata_pad_o), .SO(sdata_pad_o), .SE(scan_enable), .SI(scan_data_in));
SDFFNSRN u0_slt0_r_reg_b14_b (.CK(bit_clk_pad_i), .D(n_11436), .Q(u0_slt0_r_14), .SO(u0_slt0_r_14), .SE(scan_enable), .SI(sdata_pad_o));
SDFFNSRN u0_slt0_r_reg_b13_b (.CK(bit_clk_pad_i), .D(n_11435), .Q(u0_slt0_r_13), .SO(u0_slt0_r_13), .SE(scan_enable), .SI(u0_slt0_r_14));
SDFFNSRN u0_slt0_r_reg_b12_b (.CK(bit_clk_pad_i), .D(n_11434), .Q(u0_slt0_r_12), .SO(u0_slt0_r_12), .SE(scan_enable), .SI(u0_slt0_r_13));
SDFFNSRN u0_slt0_r_reg_b11_b (.CK(bit_clk_pad_i), .D(n_11433), .Q(u0_slt0_r_11), .SO(u0_slt0_r_11), .SE(scan_enable), .SI(u0_slt0_r_12));
SDFFNSRN u0_slt0_r_reg_b10_b (.CK(bit_clk_pad_i), .D(n_11431), .Q(u0_slt0_r_10), .SO(u0_slt0_r_10), .SE(scan_enable), .SI(u0_slt0_r_11));
SDFFNSRN u0_slt0_r_reg_b9_b (.CK(bit_clk_pad_i), .D(n_11430), .Q(u0_slt0_r_9), .SO(u0_slt0_r_9), .SE(scan_enable), .SI(u0_slt0_r_10));
SDFFNSRN u0_slt0_r_reg_b8_b (.CK(bit_clk_pad_i), .D(n_11429), .Q(u0_slt0_r_8), .SO(u0_slt0_r_8), .SE(scan_enable), .SI(u0_slt0_r_9));
SDFFNSRN u0_slt0_r_reg_b7_b (.CK(bit_clk_pad_i), .D(n_11428), .Q(u0_slt0_r_7), .SO(u0_slt0_r_7), .SE(scan_enable), .SI(u0_slt0_r_8));
SDFFNSRN u0_slt0_r_reg_b6_b (.CK(bit_clk_pad_i), .D(n_11427), .Q(u0_slt0_r_6), .SO(u0_slt0_r_6), .SE(scan_enable), .SI(u0_slt0_r_7));
SDFFNSRN u0_slt0_r_reg_b5_b (.CK(bit_clk_pad_i), .D(n_11424), .Q(u0_slt0_r_5), .SO(u0_slt0_r_5), .SE(scan_enable), .SI(u0_slt0_r_6));
SDFFNSRN u0_slt0_r_reg_b4_b (.CK(bit_clk_pad_i), .D(n_11423), .Q(u0_slt0_r_4), .SO(u0_slt0_r_4), .SE(scan_enable), .SI(u0_slt0_r_5));
SDFFNSRN u0_slt0_r_reg_b3_b (.CK(bit_clk_pad_i), .D(n_11421), .Q(u0_slt0_r_3), .SO(u0_slt0_r_3), .SE(scan_enable), .SI(u0_slt0_r_4));
SDFFNSRN u0_slt0_r_reg_b2_b (.CK(bit_clk_pad_i), .D(n_11420), .Q(u0_slt0_r_2), .SO(u0_slt0_r_2), .SE(scan_enable), .SI(u0_slt0_r_3));
SDFFNSRN u0_slt0_r_reg_b1_b (.CK(bit_clk_pad_i), .D(n_11419), .Q(u0_slt0_r_1), .SO(u0_slt0_r_1), .SE(scan_enable), .SI(u0_slt0_r_2));
SDFFNSRN u0_slt0_r_reg_b0_b (.CK(bit_clk_pad_i), .D(n_11418), .Q(u0_slt0_r), .SO(u0_slt0_r), .SE(scan_enable), .SI(u0_slt0_r_1));
SDFFNSRN u0_slt1_r_reg_b19_b (.CK(bit_clk_pad_i), .D(n_11417), .Q(u0_slt1_r_34), .SO(u0_slt1_r_34), .SE(scan_enable), .SI(u0_slt0_r));
SDFFNSRN u0_slt1_r_reg_b18_b (.CK(bit_clk_pad_i), .D(n_11416), .Q(u0_slt1_r_33), .SO(u0_slt1_r_33), .SE(scan_enable), .SI(u0_slt1_r_34));
SDFFNSRN u0_slt1_r_reg_b17_b (.CK(bit_clk_pad_i), .D(n_11414), .Q(u0_slt1_r_32), .SO(u0_slt1_r_32), .SE(scan_enable), .SI(u0_slt1_r_33));
SDFFNSRN u0_slt1_r_reg_b16_b (.CK(bit_clk_pad_i), .D(n_11413), .Q(u0_slt1_r_31), .SO(u0_slt1_r_31), .SE(scan_enable), .SI(u0_slt1_r_32));
SDFFNSRN u0_slt1_r_reg_b15_b (.CK(bit_clk_pad_i), .D(n_11411), .Q(u0_slt1_r_30), .SO(u0_slt1_r_30), .SE(scan_enable), .SI(u0_slt1_r_31));
SDFFNSRN u0_slt1_r_reg_b14_b (.CK(bit_clk_pad_i), .D(n_11410), .Q(u0_slt1_r_29), .SO(u0_slt1_r_29), .SE(scan_enable), .SI(u0_slt1_r_30));
SDFFNSRN u0_slt1_r_reg_b13_b (.CK(bit_clk_pad_i), .D(n_11409), .Q(u0_slt1_r_28), .SO(u0_slt1_r_28), .SE(scan_enable), .SI(u0_slt1_r_29));
SDFFNSRN u0_slt1_r_reg_b12_b (.CK(bit_clk_pad_i), .D(n_11408), .Q(u0_slt1_r_27), .SO(u0_slt1_r_27), .SE(scan_enable), .SI(u0_slt1_r_28));
SDFFNSRN u0_slt1_r_reg_b11_b (.CK(bit_clk_pad_i), .D(n_11406), .Q(u0_slt1_r_26), .SO(u0_slt1_r_26), .SE(scan_enable), .SI(u0_slt1_r_27));
SDFFNSRN u0_slt1_r_reg_b10_b (.CK(bit_clk_pad_i), .D(n_11404), .Q(u0_slt1_r_25), .SO(u0_slt1_r_25), .SE(scan_enable), .SI(u0_slt1_r_26));
SDFFNSRN u0_slt1_r_reg_b9_b (.CK(bit_clk_pad_i), .D(n_11403), .Q(u0_slt1_r_24), .SO(u0_slt1_r_24), .SE(scan_enable), .SI(u0_slt1_r_25));
SDFFNSRN u0_slt1_r_reg_b8_b (.CK(bit_clk_pad_i), .D(n_11401), .Q(u0_slt1_r_23), .SO(u0_slt1_r_23), .SE(scan_enable), .SI(u0_slt1_r_24));
SDFFNSRN u0_slt1_r_reg_b7_b (.CK(bit_clk_pad_i), .D(n_11400), .Q(u0_slt1_r_22), .SO(u0_slt1_r_22), .SE(scan_enable), .SI(u0_slt1_r_23));
SDFFNSRN u0_slt1_r_reg_b6_b (.CK(bit_clk_pad_i), .D(n_11399), .Q(u0_slt1_r_21), .SO(u0_slt1_r_21), .SE(scan_enable), .SI(u0_slt1_r_22));
SDFFNSRN u0_slt1_r_reg_b5_b (.CK(bit_clk_pad_i), .D(n_11397), .Q(u0_slt1_r_20), .SO(u0_slt1_r_20), .SE(scan_enable), .SI(u0_slt1_r_21));
SDFFNSRN u0_slt1_r_reg_b4_b (.CK(bit_clk_pad_i), .D(n_11396), .Q(u0_slt1_r_19), .SO(u0_slt1_r_19), .SE(scan_enable), .SI(u0_slt1_r_20));
SDFFNSRN u0_slt1_r_reg_b3_b (.CK(bit_clk_pad_i), .D(n_11394), .Q(u0_slt1_r_18), .SO(u0_slt1_r_18), .SE(scan_enable), .SI(u0_slt1_r_19));
SDFFNSRN u0_slt1_r_reg_b2_b (.CK(bit_clk_pad_i), .D(n_11393), .Q(u0_slt1_r_17), .SO(u0_slt1_r_17), .SE(scan_enable), .SI(u0_slt1_r_18));
SDFFNSRN u0_slt1_r_reg_b1_b (.CK(bit_clk_pad_i), .D(n_11392), .Q(u0_slt1_r_16), .SO(u0_slt1_r_16), .SE(scan_enable), .SI(u0_slt1_r_17));
SDFFNSRN u0_slt1_r_reg_b0_b (.CK(bit_clk_pad_i), .D(n_11391), .Q(u0_slt1_r), .SO(u0_slt1_r), .SE(scan_enable), .SI(u0_slt1_r_16));
SDFFNSRN u0_slt2_r_reg_b19_b (.CK(bit_clk_pad_i), .D(n_11390), .Q(u0_slt2_r_53), .SO(u0_slt2_r_53), .SE(scan_enable), .SI(u0_slt1_r));
SDFFNSRN u0_slt2_r_reg_b18_b (.CK(bit_clk_pad_i), .D(n_11388), .Q(u0_slt2_r_52), .SO(u0_slt2_r_52), .SE(scan_enable), .SI(u0_slt2_r_53));
SDFFNSRN u0_slt2_r_reg_b17_b (.CK(bit_clk_pad_i), .D(n_11387), .Q(u0_slt2_r_51), .SO(u0_slt2_r_51), .SE(scan_enable), .SI(u0_slt2_r_52));
SDFFNSRN u0_slt2_r_reg_b16_b (.CK(bit_clk_pad_i), .D(n_11385), .Q(u0_slt2_r_50), .SO(u0_slt2_r_50), .SE(scan_enable), .SI(u0_slt2_r_51));
SDFFNSRN u0_slt2_r_reg_b15_b (.CK(bit_clk_pad_i), .D(n_11384), .Q(u0_slt2_r_49), .SO(u0_slt2_r_49), .SE(scan_enable), .SI(u0_slt2_r_50));
SDFFNSRN u0_slt2_r_reg_b14_b (.CK(bit_clk_pad_i), .D(n_11383), .Q(u0_slt2_r_48), .SO(u0_slt2_r_48), .SE(scan_enable), .SI(u0_slt2_r_49));
SDFFNSRN u0_slt2_r_reg_b13_b (.CK(bit_clk_pad_i), .D(n_11381), .Q(u0_slt2_r_47), .SO(u0_slt2_r_47), .SE(scan_enable), .SI(u0_slt2_r_48));
SDFFNSRN u0_slt2_r_reg_b12_b (.CK(bit_clk_pad_i), .D(n_11379), .Q(u0_slt2_r_46), .SO(u0_slt2_r_46), .SE(scan_enable), .SI(u0_slt2_r_47));
SDFFNSRN u0_slt2_r_reg_b11_b (.CK(bit_clk_pad_i), .D(n_11378), .Q(u0_slt2_r_45), .SO(u0_slt2_r_45), .SE(scan_enable), .SI(u0_slt2_r_46));
SDFFNSRN u0_slt2_r_reg_b10_b (.CK(bit_clk_pad_i), .D(n_11377), .Q(u0_slt2_r_44), .SO(u0_slt2_r_44), .SE(scan_enable), .SI(u0_slt2_r_45));
SDFFNSRN u0_slt2_r_reg_b9_b (.CK(bit_clk_pad_i), .D(n_11376), .Q(u0_slt2_r_43), .SO(u0_slt2_r_43), .SE(scan_enable), .SI(u0_slt2_r_44));
SDFFNSRN u0_slt2_r_reg_b8_b (.CK(bit_clk_pad_i), .D(n_11375), .Q(u0_slt2_r_42), .SO(u0_slt2_r_42), .SE(scan_enable), .SI(u0_slt2_r_43));
SDFFNSRN u0_slt2_r_reg_b7_b (.CK(bit_clk_pad_i), .D(n_11373), .Q(u0_slt2_r_41), .SO(u0_slt2_r_41), .SE(scan_enable), .SI(u0_slt2_r_42));
SDFFNSRN u0_slt2_r_reg_b6_b (.CK(bit_clk_pad_i), .D(n_11372), .Q(u0_slt2_r_40), .SO(u0_slt2_r_40), .SE(scan_enable), .SI(u0_slt2_r_41));
SDFFNSRN u0_slt2_r_reg_b5_b (.CK(bit_clk_pad_i), .D(n_11371), .Q(u0_slt2_r_39), .SO(u0_slt2_r_39), .SE(scan_enable), .SI(u0_slt2_r_40));
SDFFNSRN u0_slt2_r_reg_b4_b (.CK(bit_clk_pad_i), .D(n_11370), .Q(u0_slt2_r_38), .SO(u0_slt2_r_38), .SE(scan_enable), .SI(u0_slt2_r_39));
SDFFNSRN u0_slt2_r_reg_b3_b (.CK(bit_clk_pad_i), .D(n_11368), .Q(u0_slt2_r_37), .SO(u0_slt2_r_37), .SE(scan_enable), .SI(u0_slt2_r_38));
SDFFNSRN u0_slt2_r_reg_b2_b (.CK(bit_clk_pad_i), .D(n_11366), .Q(u0_slt2_r_36), .SO(u0_slt2_r_36), .SE(scan_enable), .SI(u0_slt2_r_37));
SDFFNSRN u0_slt2_r_reg_b1_b (.CK(bit_clk_pad_i), .D(n_11365), .Q(u0_slt2_r_35), .SO(u0_slt2_r_35), .SE(scan_enable), .SI(u0_slt2_r_36));
SDFFNSRN u0_slt2_r_reg_b0_b (.CK(bit_clk_pad_i), .D(n_11364), .Q(u0_slt2_r), .SO(u0_slt2_r), .SE(scan_enable), .SI(u0_slt2_r_35));
SDFFNSRN u0_slt3_r_reg_b19_b (.CK(bit_clk_pad_i), .D(n_11363), .Q(u0_slt3_r_72), .SO(u0_slt3_r_72), .SE(scan_enable), .SI(u0_slt2_r));
SDFFNSRN u0_slt3_r_reg_b18_b (.CK(bit_clk_pad_i), .D(n_11361), .Q(u0_slt3_r_71), .SO(u0_slt3_r_71), .SE(scan_enable), .SI(u0_slt3_r_72));
SDFFNSRN u0_slt3_r_reg_b17_b (.CK(bit_clk_pad_i), .D(n_11360), .Q(u0_slt3_r_70), .SO(u0_slt3_r_70), .SE(scan_enable), .SI(u0_slt3_r_71));
SDFFNSRN u0_slt3_r_reg_b16_b (.CK(bit_clk_pad_i), .D(n_11358), .Q(u0_slt3_r_69), .SO(u0_slt3_r_69), .SE(scan_enable), .SI(u0_slt3_r_70));
SDFFNSRN u0_slt3_r_reg_b15_b (.CK(bit_clk_pad_i), .D(n_11356), .Q(u0_slt3_r_68), .SO(u0_slt3_r_68), .SE(scan_enable), .SI(u0_slt3_r_69));
SDFFNSRN u0_slt3_r_reg_b14_b (.CK(bit_clk_pad_i), .D(n_11355), .Q(u0_slt3_r_67), .SO(u0_slt3_r_67), .SE(scan_enable), .SI(u0_slt3_r_68));
SDFFNSRN u0_slt3_r_reg_b13_b (.CK(bit_clk_pad_i), .D(n_11354), .Q(u0_slt3_r_66), .SO(u0_slt3_r_66), .SE(scan_enable), .SI(u0_slt3_r_67));
SDFFNSRN u0_slt3_r_reg_b12_b (.CK(bit_clk_pad_i), .D(n_11353), .Q(u0_slt3_r_65), .SO(u0_slt3_r_65), .SE(scan_enable), .SI(u0_slt3_r_66));
SDFFNSRN u0_slt3_r_reg_b11_b (.CK(bit_clk_pad_i), .D(n_11352), .Q(u0_slt3_r_64), .SO(u0_slt3_r_64), .SE(scan_enable), .SI(u0_slt3_r_65));
SDFFNSRN u0_slt3_r_reg_b10_b (.CK(bit_clk_pad_i), .D(n_11351), .Q(u0_slt3_r_63), .SO(u0_slt3_r_63), .SE(scan_enable), .SI(u0_slt3_r_64));
SDFFNSRN u0_slt3_r_reg_b9_b (.CK(bit_clk_pad_i), .D(n_11349), .Q(u0_slt3_r_62), .SO(u0_slt3_r_62), .SE(scan_enable), .SI(u0_slt3_r_63));
SDFFNSRN u0_slt3_r_reg_b8_b (.CK(bit_clk_pad_i), .D(n_11348), .Q(u0_slt3_r_61), .SO(u0_slt3_r_61), .SE(scan_enable), .SI(u0_slt3_r_62));
SDFFNSRN u0_slt3_r_reg_b7_b (.CK(bit_clk_pad_i), .D(n_11347), .Q(u0_slt3_r_60), .SO(u0_slt3_r_60), .SE(scan_enable), .SI(u0_slt3_r_61));
SDFFNSRN u0_slt3_r_reg_b6_b (.CK(bit_clk_pad_i), .D(n_11346), .Q(u0_slt3_r_59), .SO(u0_slt3_r_59), .SE(scan_enable), .SI(u0_slt3_r_60));
SDFFNSRN u0_slt3_r_reg_b5_b (.CK(bit_clk_pad_i), .D(n_11344), .Q(u0_slt3_r_58), .SO(u0_slt3_r_58), .SE(scan_enable), .SI(u0_slt3_r_59));
SDFFNSRN u0_slt3_r_reg_b4_b (.CK(bit_clk_pad_i), .D(n_11342), .Q(u0_slt3_r_57), .SO(u0_slt3_r_57), .SE(scan_enable), .SI(u0_slt3_r_58));
SDFFNSRN u0_slt3_r_reg_b3_b (.CK(bit_clk_pad_i), .D(n_11341), .Q(u0_slt3_r_56), .SO(u0_slt3_r_56), .SE(scan_enable), .SI(u0_slt3_r_57));
SDFFNSRN u0_slt3_r_reg_b2_b (.CK(bit_clk_pad_i), .D(n_11339), .Q(u0_slt3_r_55), .SO(u0_slt3_r_55), .SE(scan_enable), .SI(u0_slt3_r_56));
SDFFNSRN u0_slt3_r_reg_b1_b (.CK(bit_clk_pad_i), .D(n_11338), .Q(u0_slt3_r_54), .SO(u0_slt3_r_54), .SE(scan_enable), .SI(u0_slt3_r_55));
SDFFNSRN u0_slt3_r_reg_b0_b (.CK(bit_clk_pad_i), .D(n_11336), .Q(u0_slt3_r), .SO(u0_slt3_r), .SE(scan_enable), .SI(u0_slt3_r_54));
SDFFNSRN u0_slt4_r_reg_b19_b (.CK(bit_clk_pad_i), .D(n_11334), .Q(u0_slt4_r_91), .SO(u0_slt4_r_91), .SE(scan_enable), .SI(u0_slt3_r));
SDFFNSRN u0_slt4_r_reg_b18_b (.CK(bit_clk_pad_i), .D(n_11333), .Q(u0_slt4_r_90), .SO(u0_slt4_r_90), .SE(scan_enable), .SI(u0_slt4_r_91));
SDFFNSRN u0_slt4_r_reg_b17_b (.CK(bit_clk_pad_i), .D(n_11332), .Q(u0_slt4_r_89), .SO(u0_slt4_r_89), .SE(scan_enable), .SI(u0_slt4_r_90));
SDFFNSRN u0_slt4_r_reg_b16_b (.CK(bit_clk_pad_i), .D(n_11330), .Q(u0_slt4_r_88), .SO(u0_slt4_r_88), .SE(scan_enable), .SI(u0_slt4_r_89));
SDFFNSRN u0_slt4_r_reg_b15_b (.CK(bit_clk_pad_i), .D(n_11329), .Q(u0_slt4_r_87), .SO(u0_slt4_r_87), .SE(scan_enable), .SI(u0_slt4_r_88));
SDFFNSRN u0_slt4_r_reg_b14_b (.CK(bit_clk_pad_i), .D(n_11328), .Q(u0_slt4_r_86), .SO(u0_slt4_r_86), .SE(scan_enable), .SI(u0_slt4_r_87));
SDFFNSRN u0_slt4_r_reg_b13_b (.CK(bit_clk_pad_i), .D(n_11327), .Q(u0_slt4_r_85), .SO(u0_slt4_r_85), .SE(scan_enable), .SI(u0_slt4_r_86));
SDFFNSRN u0_slt4_r_reg_b12_b (.CK(bit_clk_pad_i), .D(n_11326), .Q(u0_slt4_r_84), .SO(u0_slt4_r_84), .SE(scan_enable), .SI(u0_slt4_r_85));
SDFFNSRN u0_slt4_r_reg_b11_b (.CK(bit_clk_pad_i), .D(n_11324), .Q(u0_slt4_r_83), .SO(u0_slt4_r_83), .SE(scan_enable), .SI(u0_slt4_r_84));
SDFFNSRN u0_slt4_r_reg_b10_b (.CK(bit_clk_pad_i), .D(n_11323), .Q(u0_slt4_r_82), .SO(u0_slt4_r_82), .SE(scan_enable), .SI(u0_slt4_r_83));
SDFFNSRN u0_slt4_r_reg_b9_b (.CK(bit_clk_pad_i), .D(n_11321), .Q(u0_slt4_r_81), .SO(u0_slt4_r_81), .SE(scan_enable), .SI(u0_slt4_r_82));
SDFFNSRN u0_slt4_r_reg_b8_b (.CK(bit_clk_pad_i), .D(n_11320), .Q(u0_slt4_r_80), .SO(u0_slt4_r_80), .SE(scan_enable), .SI(u0_slt4_r_81));
SDFFNSRN u0_slt4_r_reg_b7_b (.CK(bit_clk_pad_i), .D(n_11318), .Q(u0_slt4_r_79), .SO(u0_slt4_r_79), .SE(scan_enable), .SI(u0_slt4_r_80));
SDFFNSRN u0_slt4_r_reg_b6_b (.CK(bit_clk_pad_i), .D(n_11317), .Q(u0_slt4_r_78), .SO(u0_slt4_r_78), .SE(scan_enable), .SI(u0_slt4_r_79));
SDFFNSRN u0_slt4_r_reg_b5_b (.CK(bit_clk_pad_i), .D(n_11315), .Q(u0_slt4_r_77), .SO(u0_slt4_r_77), .SE(scan_enable), .SI(u0_slt4_r_78));
SDFFNSRN u0_slt4_r_reg_b4_b (.CK(bit_clk_pad_i), .D(n_11314), .Q(u0_slt4_r_76), .SO(u0_slt4_r_76), .SE(scan_enable), .SI(u0_slt4_r_77));
SDFFNSRN u0_slt4_r_reg_b3_b (.CK(bit_clk_pad_i), .D(n_11313), .Q(u0_slt4_r_75), .SO(u0_slt4_r_75), .SE(scan_enable), .SI(u0_slt4_r_76));
SDFFNSRN u0_slt4_r_reg_b2_b (.CK(bit_clk_pad_i), .D(n_11312), .Q(u0_slt4_r_74), .SO(u0_slt4_r_74), .SE(scan_enable), .SI(u0_slt4_r_75));
SDFFNSRN u0_slt4_r_reg_b1_b (.CK(bit_clk_pad_i), .D(n_11311), .Q(u0_slt4_r_73), .SO(u0_slt4_r_73), .SE(scan_enable), .SI(u0_slt4_r_74));
SDFFNSRN u0_slt4_r_reg_b0_b (.CK(bit_clk_pad_i), .D(n_11310), .Q(u0_slt4_r), .SO(u0_slt4_r), .SE(scan_enable), .SI(u0_slt4_r_73));
SDFFNSRN u0_slt5_r_reg_b19_b (.CK(bit_clk_pad_i), .D(n_11308), .Q(u0_slt5_r_110), .SO(u0_slt5_r_110), .SE(scan_enable), .SI(u0_slt4_r));
SDFFNSRN u0_slt5_r_reg_b18_b (.CK(bit_clk_pad_i), .D(n_11307), .Q(u0_slt5_r_109), .SO(u0_slt5_r_109), .SE(scan_enable), .SI(u0_slt5_r_110));
SDFFNSRN u0_slt5_r_reg_b17_b (.CK(bit_clk_pad_i), .D(n_11306), .Q(u0_slt5_r_108), .SO(u0_slt5_r_108), .SE(scan_enable), .SI(u0_slt5_r_109));
SDFFNSRN u0_slt5_r_reg_b16_b (.CK(bit_clk_pad_i), .D(n_11305), .Q(u0_slt5_r_107), .SO(u0_slt5_r_107), .SE(scan_enable), .SI(u0_slt5_r_108));
SDFFNSRN u0_slt5_r_reg_b15_b (.CK(bit_clk_pad_i), .D(n_11304), .Q(u0_slt5_r_106), .SO(u0_slt5_r_106), .SE(scan_enable), .SI(u0_slt5_r_107));
SDFFNSRN u0_slt5_r_reg_b14_b (.CK(bit_clk_pad_i), .D(n_11303), .Q(u0_slt5_r_105), .SO(u0_slt5_r_105), .SE(scan_enable), .SI(u0_slt5_r_106));
SDFFNSRN u0_slt5_r_reg_b13_b (.CK(bit_clk_pad_i), .D(n_11302), .Q(u0_slt5_r_104), .SO(u0_slt5_r_104), .SE(scan_enable), .SI(u0_slt5_r_105));
SDFFNSRN u0_slt5_r_reg_b12_b (.CK(bit_clk_pad_i), .D(n_11301), .Q(u0_slt5_r_103), .SO(u0_slt5_r_103), .SE(scan_enable), .SI(u0_slt5_r_104));
SDFFNSRN u0_slt5_r_reg_b11_b (.CK(bit_clk_pad_i), .D(n_11300), .Q(u0_slt5_r_102), .SO(u0_slt5_r_102), .SE(scan_enable), .SI(u0_slt5_r_103));
SDFFNSRN u0_slt5_r_reg_b10_b (.CK(bit_clk_pad_i), .D(n_11299), .Q(u0_slt5_r_101), .SO(u0_slt5_r_101), .SE(scan_enable), .SI(u0_slt5_r_102));
SDFFNSRN u0_slt5_r_reg_b9_b (.CK(bit_clk_pad_i), .D(n_11298), .Q(u0_slt5_r_100), .SO(u0_slt5_r_100), .SE(scan_enable), .SI(u0_slt5_r_101));
SDFFNSRN u0_slt5_r_reg_b8_b (.CK(bit_clk_pad_i), .D(n_11297), .Q(u0_slt5_r_99), .SO(u0_slt5_r_99), .SE(scan_enable), .SI(u0_slt5_r_100));
SDFFNSRN u0_slt5_r_reg_b7_b (.CK(bit_clk_pad_i), .D(n_11296), .Q(u0_slt5_r_98), .SO(u0_slt5_r_98), .SE(scan_enable), .SI(u0_slt5_r_99));
SDFFNSRN u0_slt5_r_reg_b6_b (.CK(bit_clk_pad_i), .D(n_11295), .Q(u0_slt5_r_97), .SO(u0_slt5_r_97), .SE(scan_enable), .SI(u0_slt5_r_98));
SDFFNSRN u0_slt5_r_reg_b5_b (.CK(bit_clk_pad_i), .D(n_11294), .Q(u0_slt5_r_96), .SO(u0_slt5_r_96), .SE(scan_enable), .SI(u0_slt5_r_97));
SDFFNSRN u0_slt5_r_reg_b4_b (.CK(bit_clk_pad_i), .D(n_11293), .Q(u0_slt5_r_95), .SO(u0_slt5_r_95), .SE(scan_enable), .SI(u0_slt5_r_96));
SDFFNSRN u0_slt5_r_reg_b3_b (.CK(bit_clk_pad_i), .D(n_11292), .Q(u0_slt5_r_94), .SO(u0_slt5_r_94), .SE(scan_enable), .SI(u0_slt5_r_95));
SDFFNSRN u0_slt5_r_reg_b2_b (.CK(bit_clk_pad_i), .D(n_11291), .Q(u0_slt5_r_93), .SO(u0_slt5_r_93), .SE(scan_enable), .SI(u0_slt5_r_94));
SDFFNSRN u0_slt5_r_reg_b1_b (.CK(bit_clk_pad_i), .D(n_11290), .Q(u0_slt5_r_92), .SO(u0_slt5_r_92), .SE(scan_enable), .SI(u0_slt5_r_93));
SDFFNSRN u0_slt5_r_reg_b0_b (.CK(bit_clk_pad_i), .D(n_11289), .Q(u0_slt5_r), .SO(u0_slt5_r), .SE(scan_enable), .SI(u0_slt5_r_92));
SDFFNSRN u0_slt6_r_reg_b19_b (.CK(bit_clk_pad_i), .D(n_11288), .Q(u0_slt6_r_129), .SO(u0_slt6_r_129), .SE(scan_enable), .SI(u0_slt5_r));
SDFFNSRN u0_slt6_r_reg_b18_b (.CK(bit_clk_pad_i), .D(n_11287), .Q(u0_slt6_r_128), .SO(u0_slt6_r_128), .SE(scan_enable), .SI(u0_slt6_r_129));
SDFFNSRN u0_slt6_r_reg_b17_b (.CK(bit_clk_pad_i), .D(n_11286), .Q(u0_slt6_r_127), .SO(u0_slt6_r_127), .SE(scan_enable), .SI(u0_slt6_r_128));
SDFFNSRN u0_slt6_r_reg_b16_b (.CK(bit_clk_pad_i), .D(n_11284), .Q(u0_slt6_r_126), .SO(u0_slt6_r_126), .SE(scan_enable), .SI(u0_slt6_r_127));
SDFFNSRN u0_slt6_r_reg_b15_b (.CK(bit_clk_pad_i), .D(n_11283), .Q(u0_slt6_r_125), .SO(u0_slt6_r_125), .SE(scan_enable), .SI(u0_slt6_r_126));
SDFFNSRN u0_slt6_r_reg_b14_b (.CK(bit_clk_pad_i), .D(n_11281), .Q(u0_slt6_r_124), .SO(u0_slt6_r_124), .SE(scan_enable), .SI(u0_slt6_r_125));
SDFFNSRN u0_slt6_r_reg_b13_b (.CK(bit_clk_pad_i), .D(n_11280), .Q(u0_slt6_r_123), .SO(u0_slt6_r_123), .SE(scan_enable), .SI(u0_slt6_r_124));
SDFFNSRN u0_slt6_r_reg_b12_b (.CK(bit_clk_pad_i), .D(n_11279), .Q(u0_slt6_r_122), .SO(u0_slt6_r_122), .SE(scan_enable), .SI(u0_slt6_r_123));
SDFFNSRN u0_slt6_r_reg_b11_b (.CK(bit_clk_pad_i), .D(n_11278), .Q(u0_slt6_r_121), .SO(u0_slt6_r_121), .SE(scan_enable), .SI(u0_slt6_r_122));
SDFFNSRN u0_slt6_r_reg_b10_b (.CK(bit_clk_pad_i), .D(n_11276), .Q(u0_slt6_r_120), .SO(u0_slt6_r_120), .SE(scan_enable), .SI(u0_slt6_r_121));
SDFFNSRN u0_slt6_r_reg_b9_b (.CK(bit_clk_pad_i), .D(n_11274), .Q(u0_slt6_r_119), .SO(u0_slt6_r_119), .SE(scan_enable), .SI(u0_slt6_r_120));
SDFFNSRN u0_slt6_r_reg_b8_b (.CK(bit_clk_pad_i), .D(n_11273), .Q(u0_slt6_r_118), .SO(u0_slt6_r_118), .SE(scan_enable), .SI(u0_slt6_r_119));
SDFFNSRN u0_slt6_r_reg_b7_b (.CK(bit_clk_pad_i), .D(n_11272), .Q(u0_slt6_r_117), .SO(u0_slt6_r_117), .SE(scan_enable), .SI(u0_slt6_r_118));
SDFFNSRN u0_slt6_r_reg_b6_b (.CK(bit_clk_pad_i), .D(n_11270), .Q(u0_slt6_r_116), .SO(u0_slt6_r_116), .SE(scan_enable), .SI(u0_slt6_r_117));
SDFFNSRN u0_slt6_r_reg_b5_b (.CK(bit_clk_pad_i), .D(n_11269), .Q(u0_slt6_r_115), .SO(u0_slt6_r_115), .SE(scan_enable), .SI(u0_slt6_r_116));
SDFFNSRN u0_slt6_r_reg_b4_b (.CK(bit_clk_pad_i), .D(n_11268), .Q(u0_slt6_r_114), .SO(u0_slt6_r_114), .SE(scan_enable), .SI(u0_slt6_r_115));
SDFFNSRN u0_slt6_r_reg_b3_b (.CK(bit_clk_pad_i), .D(n_11267), .Q(u0_slt6_r_113), .SO(u0_slt6_r_113), .SE(scan_enable), .SI(u0_slt6_r_114));
SDFFNSRN u0_slt6_r_reg_b2_b (.CK(bit_clk_pad_i), .D(n_11266), .Q(u0_slt6_r_112), .SO(u0_slt6_r_112), .SE(scan_enable), .SI(u0_slt6_r_113));
SDFFNSRN u0_slt6_r_reg_b1_b (.CK(bit_clk_pad_i), .D(n_11264), .Q(u0_slt6_r_111), .SO(u0_slt6_r_111), .SE(scan_enable), .SI(u0_slt6_r_112));
SDFFNSRN u0_slt6_r_reg_b0_b (.CK(bit_clk_pad_i), .D(n_11263), .Q(u0_slt6_r), .SO(u0_slt6_r), .SE(scan_enable), .SI(u0_slt6_r_111));
SDFFNSRN u0_slt7_r_reg_b19_b (.CK(bit_clk_pad_i), .D(n_11262), .Q(u0_slt7_r_148), .SO(u0_slt7_r_148), .SE(scan_enable), .SI(u0_slt6_r));
SDFFNSRN u0_slt7_r_reg_b18_b (.CK(bit_clk_pad_i), .D(n_11260), .Q(u0_slt7_r_147), .SO(u0_slt7_r_147), .SE(scan_enable), .SI(u0_slt7_r_148));
SDFFNSRN u0_slt7_r_reg_b17_b (.CK(bit_clk_pad_i), .D(n_11258), .Q(u0_slt7_r_146), .SO(u0_slt7_r_146), .SE(scan_enable), .SI(u0_slt7_r_147));
SDFFNSRN u0_slt7_r_reg_b16_b (.CK(bit_clk_pad_i), .D(n_11257), .Q(u0_slt7_r_145), .SO(u0_slt7_r_145), .SE(scan_enable), .SI(u0_slt7_r_146));
SDFFNSRN u0_slt7_r_reg_b15_b (.CK(bit_clk_pad_i), .D(n_11256), .Q(u0_slt7_r_144), .SO(u0_slt7_r_144), .SE(scan_enable), .SI(u0_slt7_r_145));
SDFFNSRN u0_slt7_r_reg_b14_b (.CK(bit_clk_pad_i), .D(n_11255), .Q(u0_slt7_r_143), .SO(u0_slt7_r_143), .SE(scan_enable), .SI(u0_slt7_r_144));
SDFFNSRN u0_slt7_r_reg_b13_b (.CK(bit_clk_pad_i), .D(n_11254), .Q(u0_slt7_r_142), .SO(u0_slt7_r_142), .SE(scan_enable), .SI(u0_slt7_r_143));
SDFFNSRN u0_slt7_r_reg_b12_b (.CK(bit_clk_pad_i), .D(n_11253), .Q(u0_slt7_r_141), .SO(u0_slt7_r_141), .SE(scan_enable), .SI(u0_slt7_r_142));
SDFFNSRN u0_slt7_r_reg_b11_b (.CK(bit_clk_pad_i), .D(n_11252), .Q(u0_slt7_r_140), .SO(u0_slt7_r_140), .SE(scan_enable), .SI(u0_slt7_r_141));
SDFFNSRN u0_slt7_r_reg_b10_b (.CK(bit_clk_pad_i), .D(n_11251), .Q(u0_slt7_r_139), .SO(u0_slt7_r_139), .SE(scan_enable), .SI(u0_slt7_r_140));
SDFFNSRN u0_slt7_r_reg_b9_b (.CK(bit_clk_pad_i), .D(n_11250), .Q(u0_slt7_r_138), .SO(u0_slt7_r_138), .SE(scan_enable), .SI(u0_slt7_r_139));
SDFFNSRN u0_slt7_r_reg_b8_b (.CK(bit_clk_pad_i), .D(n_11249), .Q(u0_slt7_r_137), .SO(u0_slt7_r_137), .SE(scan_enable), .SI(u0_slt7_r_138));
SDFFNSRN u0_slt7_r_reg_b7_b (.CK(bit_clk_pad_i), .D(n_11248), .Q(u0_slt7_r_136), .SO(u0_slt7_r_136), .SE(scan_enable), .SI(u0_slt7_r_137));
SDFFNSRN u0_slt7_r_reg_b6_b (.CK(bit_clk_pad_i), .D(n_11247), .Q(u0_slt7_r_135), .SO(u0_slt7_r_135), .SE(scan_enable), .SI(u0_slt7_r_136));
SDFFNSRN u0_slt7_r_reg_b5_b (.CK(bit_clk_pad_i), .D(n_11246), .Q(u0_slt7_r_134), .SO(u0_slt7_r_134), .SE(scan_enable), .SI(u0_slt7_r_135));
SDFFNSRN u0_slt7_r_reg_b4_b (.CK(bit_clk_pad_i), .D(n_11245), .Q(u0_slt7_r_133), .SO(u0_slt7_r_133), .SE(scan_enable), .SI(u0_slt7_r_134));
SDFFNSRN u0_slt7_r_reg_b3_b (.CK(bit_clk_pad_i), .D(n_11244), .Q(u0_slt7_r_132), .SO(u0_slt7_r_132), .SE(scan_enable), .SI(u0_slt7_r_133));
SDFFNSRN u0_slt7_r_reg_b2_b (.CK(bit_clk_pad_i), .D(n_11243), .Q(u0_slt7_r_131), .SO(u0_slt7_r_131), .SE(scan_enable), .SI(u0_slt7_r_132));
SDFFNSRN u0_slt7_r_reg_b1_b (.CK(bit_clk_pad_i), .D(n_11242), .Q(u0_slt7_r_130), .SO(u0_slt7_r_130), .SE(scan_enable), .SI(u0_slt7_r_131));
SDFFNSRN u0_slt7_r_reg_b0_b (.CK(bit_clk_pad_i), .D(n_11241), .Q(u0_slt7_r), .SO(u0_slt7_r), .SE(scan_enable), .SI(u0_slt7_r_130));
SDFFNSRN u0_slt8_r_reg_b19_b (.CK(bit_clk_pad_i), .D(n_11240), .Q(u0_slt8_r_167), .SO(u0_slt8_r_167), .SE(scan_enable), .SI(u0_slt7_r));
SDFFNSRN u0_slt8_r_reg_b18_b (.CK(bit_clk_pad_i), .D(n_11239), .Q(u0_slt8_r_166), .SO(u0_slt8_r_166), .SE(scan_enable), .SI(u0_slt8_r_167));
SDFFNSRN u0_slt8_r_reg_b17_b (.CK(bit_clk_pad_i), .D(n_11238), .Q(u0_slt8_r_165), .SO(u0_slt8_r_165), .SE(scan_enable), .SI(u0_slt8_r_166));
SDFFNSRN u0_slt8_r_reg_b16_b (.CK(bit_clk_pad_i), .D(n_11237), .Q(u0_slt8_r_164), .SO(u0_slt8_r_164), .SE(scan_enable), .SI(u0_slt8_r_165));
SDFFNSRN u0_slt8_r_reg_b15_b (.CK(bit_clk_pad_i), .D(n_11236), .Q(u0_slt8_r_163), .SO(u0_slt8_r_163), .SE(scan_enable), .SI(u0_slt8_r_164));
SDFFNSRN u0_slt8_r_reg_b14_b (.CK(bit_clk_pad_i), .D(n_11235), .Q(u0_slt8_r_162), .SO(u0_slt8_r_162), .SE(scan_enable), .SI(u0_slt8_r_163));
SDFFNSRN u0_slt8_r_reg_b13_b (.CK(bit_clk_pad_i), .D(n_11234), .Q(u0_slt8_r_161), .SO(u0_slt8_r_161), .SE(scan_enable), .SI(u0_slt8_r_162));
SDFFNSRN u0_slt8_r_reg_b12_b (.CK(bit_clk_pad_i), .D(n_11233), .Q(u0_slt8_r_160), .SO(u0_slt8_r_160), .SE(scan_enable), .SI(u0_slt8_r_161));
SDFFNSRN u0_slt8_r_reg_b11_b (.CK(bit_clk_pad_i), .D(n_11232), .Q(u0_slt8_r_159), .SO(u0_slt8_r_159), .SE(scan_enable), .SI(u0_slt8_r_160));
SDFFNSRN u0_slt8_r_reg_b10_b (.CK(bit_clk_pad_i), .D(n_11231), .Q(u0_slt8_r_158), .SO(u0_slt8_r_158), .SE(scan_enable), .SI(u0_slt8_r_159));
SDFFNSRN u0_slt8_r_reg_b9_b (.CK(bit_clk_pad_i), .D(n_11230), .Q(u0_slt8_r_157), .SO(u0_slt8_r_157), .SE(scan_enable), .SI(u0_slt8_r_158));
SDFFNSRN u0_slt8_r_reg_b8_b (.CK(bit_clk_pad_i), .D(n_11228), .Q(u0_slt8_r_156), .SO(u0_slt8_r_156), .SE(scan_enable), .SI(u0_slt8_r_157));
SDFFNSRN u0_slt8_r_reg_b7_b (.CK(bit_clk_pad_i), .D(n_11227), .Q(u0_slt8_r_155), .SO(u0_slt8_r_155), .SE(scan_enable), .SI(u0_slt8_r_156));
SDFFNSRN u0_slt8_r_reg_b6_b (.CK(bit_clk_pad_i), .D(n_11225), .Q(u0_slt8_r_154), .SO(u0_slt8_r_154), .SE(scan_enable), .SI(u0_slt8_r_155));
SDFFNSRN u0_slt8_r_reg_b5_b (.CK(bit_clk_pad_i), .D(n_11224), .Q(u0_slt8_r_153), .SO(u0_slt8_r_153), .SE(scan_enable), .SI(u0_slt8_r_154));
SDFFNSRN u0_slt8_r_reg_b4_b (.CK(bit_clk_pad_i), .D(n_11223), .Q(u0_slt8_r_152), .SO(u0_slt8_r_152), .SE(scan_enable), .SI(u0_slt8_r_153));
SDFFNSRN u0_slt8_r_reg_b3_b (.CK(bit_clk_pad_i), .D(n_11221), .Q(u0_slt8_r_151), .SO(u0_slt8_r_151), .SE(scan_enable), .SI(u0_slt8_r_152));
SDFFNSRN u0_slt8_r_reg_b2_b (.CK(bit_clk_pad_i), .D(n_11220), .Q(u0_slt8_r_150), .SO(u0_slt8_r_150), .SE(scan_enable), .SI(u0_slt8_r_151));
SDFFNSRN u0_slt8_r_reg_b1_b (.CK(bit_clk_pad_i), .D(n_11219), .Q(u0_slt8_r_149), .SO(u0_slt8_r_149), .SE(scan_enable), .SI(u0_slt8_r_150));
SDFFNSRN u0_slt8_r_reg_b0_b (.CK(bit_clk_pad_i), .D(n_11218), .Q(u0_slt8_r), .SO(u0_slt8_r), .SE(scan_enable), .SI(u0_slt8_r_149));
SDFFNSRN u0_slt9_r_reg_b19_b (.CK(bit_clk_pad_i), .D(n_11217), .Q(u0_slt9_r_186), .SO(u0_slt9_r_186), .SE(scan_enable), .SI(u0_slt8_r));
SDFFNSRN u0_slt9_r_reg_b18_b (.CK(bit_clk_pad_i), .D(n_11216), .Q(u0_slt9_r_185), .SO(u0_slt9_r_185), .SE(scan_enable), .SI(u0_slt9_r_186));
SDFFNSRN u0_slt9_r_reg_b17_b (.CK(bit_clk_pad_i), .D(n_11215), .Q(u0_slt9_r_184), .SO(u0_slt9_r_184), .SE(scan_enable), .SI(u0_slt9_r_185));
SDFFNSRN u0_slt9_r_reg_b16_b (.CK(bit_clk_pad_i), .D(n_11214), .Q(u0_slt9_r_183), .SO(u0_slt9_r_183), .SE(scan_enable), .SI(u0_slt9_r_184));
SDFFNSRN u0_slt9_r_reg_b15_b (.CK(bit_clk_pad_i), .D(n_11213), .Q(u0_slt9_r_182), .SO(u0_slt9_r_182), .SE(scan_enable), .SI(u0_slt9_r_183));
SDFFNSRN u0_slt9_r_reg_b14_b (.CK(bit_clk_pad_i), .D(n_11212), .Q(u0_slt9_r_181), .SO(u0_slt9_r_181), .SE(scan_enable), .SI(u0_slt9_r_182));
SDFFNSRN u0_slt9_r_reg_b13_b (.CK(bit_clk_pad_i), .D(n_11211), .Q(u0_slt9_r_180), .SO(u0_slt9_r_180), .SE(scan_enable), .SI(u0_slt9_r_181));
SDFFNSRN u0_slt9_r_reg_b12_b (.CK(bit_clk_pad_i), .D(n_11210), .Q(u0_slt9_r_179), .SO(u0_slt9_r_179), .SE(scan_enable), .SI(u0_slt9_r_180));
SDFFNSRN u0_slt9_r_reg_b11_b (.CK(bit_clk_pad_i), .D(n_11209), .Q(u0_slt9_r_178), .SO(u0_slt9_r_178), .SE(scan_enable), .SI(u0_slt9_r_179));
SDFFNSRN u0_slt9_r_reg_b10_b (.CK(bit_clk_pad_i), .D(n_11207), .Q(u0_slt9_r_177), .SO(u0_slt9_r_177), .SE(scan_enable), .SI(u0_slt9_r_178));
SDFFNSRN u0_slt9_r_reg_b9_b (.CK(bit_clk_pad_i), .D(n_11206), .Q(u0_slt9_r_176), .SO(u0_slt9_r_176), .SE(scan_enable), .SI(u0_slt9_r_177));
SDFFNSRN u0_slt9_r_reg_b8_b (.CK(bit_clk_pad_i), .D(n_11205), .Q(u0_slt9_r_175), .SO(u0_slt9_r_175), .SE(scan_enable), .SI(u0_slt9_r_176));
SDFFNSRN u0_slt9_r_reg_b7_b (.CK(bit_clk_pad_i), .D(n_11204), .Q(u0_slt9_r_174), .SO(u0_slt9_r_174), .SE(scan_enable), .SI(u0_slt9_r_175));
SDFFNSRN u0_slt9_r_reg_b6_b (.CK(bit_clk_pad_i), .D(n_11203), .Q(u0_slt9_r_173), .SO(u0_slt9_r_173), .SE(scan_enable), .SI(u0_slt9_r_174));
SDFFNSRN u1_slt2_reg_b19_b (.CK(bit_clk_pad_i), .D(n_11202), .Q(in_slt_845), .SO(in_slt_845), .SE(scan_enable), .SI(u0_slt9_r_173));
SDFFNSRN u1_slt3_reg_b19_b (.CK(bit_clk_pad_i), .D(n_11201), .Q(in_slt_415), .SO(in_slt_415), .SE(scan_enable), .SI(in_slt_845));
SDFFNSRN u1_slt4_reg_b19_b (.CK(bit_clk_pad_i), .D(n_11200), .Q(in_slt_437), .SO(in_slt_437), .SE(scan_enable), .SI(in_slt_415));
SDFFNSRN u1_slt6_reg_b19_b (.CK(bit_clk_pad_i), .D(n_11199), .Q(in_slt_459), .SO(in_slt_459), .SE(scan_enable), .SI(in_slt_437));
SDFFNSRN u1_slt2_reg_b18_b (.CK(bit_clk_pad_i), .D(n_11198), .Q(in_slt_844), .SO(in_slt_844), .SE(scan_enable), .SI(in_slt_459));
SDFFNSRN u1_slt3_reg_b18_b (.CK(bit_clk_pad_i), .D(n_11197), .Q(in_slt_414), .SO(in_slt_414), .SE(scan_enable), .SI(in_slt_844));
SDFFNSRN u1_slt4_reg_b18_b (.CK(bit_clk_pad_i), .D(n_11196), .Q(in_slt_436), .SO(in_slt_436), .SE(scan_enable), .SI(in_slt_414));
SDFFNSRN u1_slt6_reg_b18_b (.CK(bit_clk_pad_i), .D(n_11195), .Q(in_slt_458), .SO(in_slt_458), .SE(scan_enable), .SI(in_slt_436));
SDFFNSRN u0_slt9_r_reg_b5_b (.CK(bit_clk_pad_i), .D(n_11188), .Q(u0_slt9_r_172), .SO(u0_slt9_r_172), .SE(scan_enable), .SI(in_slt_458));
SDFFNSRN u1_slt2_reg_b17_b (.CK(bit_clk_pad_i), .D(n_11187), .Q(in_slt_843), .SO(in_slt_843), .SE(scan_enable), .SI(u0_slt9_r_172));
SDFFNSRN u1_slt3_reg_b17_b (.CK(bit_clk_pad_i), .D(n_11186), .Q(in_slt_413), .SO(in_slt_413), .SE(scan_enable), .SI(in_slt_843));
SDFFNSRN u1_slt4_reg_b17_b (.CK(bit_clk_pad_i), .D(n_11185), .Q(in_slt_435), .SO(in_slt_435), .SE(scan_enable), .SI(in_slt_413));
SDFFNSRN u1_slt6_reg_b17_b (.CK(bit_clk_pad_i), .D(n_11184), .Q(in_slt_457), .SO(in_slt_457), .SE(scan_enable), .SI(in_slt_435));
SDFFNSRN u1_sr_reg_b19_b (.CK(bit_clk_pad_i), .D(u1_sr_134), .Q(u1_sr_135), .SO(u1_sr_135), .SE(scan_enable), .SI(in_slt_457));
SDFFNSRN u1_slt2_reg_b16_b (.CK(bit_clk_pad_i), .D(n_11169), .Q(in_slt_842), .SO(in_slt_842), .SE(scan_enable), .SI(u1_sr_135));
SDFFNSRN u1_slt3_reg_b16_b (.CK(bit_clk_pad_i), .D(n_11168), .Q(in_slt_412), .SO(in_slt_412), .SE(scan_enable), .SI(in_slt_842));
SDFFNSRN u1_slt4_reg_b16_b (.CK(bit_clk_pad_i), .D(n_11167), .Q(in_slt_434), .SO(in_slt_434), .SE(scan_enable), .SI(in_slt_412));
SDFFNSRN u1_slt6_reg_b16_b (.CK(bit_clk_pad_i), .D(n_11166), .Q(in_slt_456), .SO(in_slt_456), .SE(scan_enable), .SI(in_slt_434));
SDFFNSRN u1_sr_reg_b18_b (.CK(bit_clk_pad_i), .D(u1_sr_133), .Q(u1_sr_134), .SO(u1_sr_134), .SE(scan_enable), .SI(in_slt_456));
SDFFNSRN u1_slt3_reg_b15_b (.CK(bit_clk_pad_i), .D(n_11116), .Q(in_slt_411), .SO(in_slt_411), .SE(scan_enable), .SI(u1_sr_134));
SDFFNSRN u1_slt0_reg_b15_b (.CK(bit_clk_pad_i), .D(n_11118), .Q(in_slt_742), .SO(in_slt_742), .SE(scan_enable), .SI(in_slt_411));
SDFFNSRN u1_slt6_reg_b15_b (.CK(bit_clk_pad_i), .D(n_11114), .Q(in_slt_455), .SO(in_slt_455), .SE(scan_enable), .SI(in_slt_742));
SDFFNSRN u1_slt2_reg_b15_b (.CK(bit_clk_pad_i), .D(n_11117), .Q(in_slt_841), .SO(in_slt_841), .SE(scan_enable), .SI(in_slt_455));
SDFFNSRN u1_slt4_reg_b15_b (.CK(bit_clk_pad_i), .D(n_11115), .Q(in_slt_433), .SO(in_slt_433), .SE(scan_enable), .SI(in_slt_841));
SDFFNSRN u0_slt9_r_reg_b4_b (.CK(bit_clk_pad_i), .D(n_11010), .Q(u0_slt9_r_171), .SO(u0_slt9_r_171), .SE(scan_enable), .SI(in_slt_433));
SDFFNSRN u1_sr_reg_b17_b (.CK(bit_clk_pad_i), .D(u1_sr_132), .Q(u1_sr_133), .SO(u1_sr_133), .SE(scan_enable), .SI(u0_slt9_r_171));
SDFFNSRN u1_slt3_reg_b14_b (.CK(bit_clk_pad_i), .D(n_10961), .Q(in_slt_410), .SO(in_slt_410), .SE(scan_enable), .SI(u1_sr_133));
SDFFNSRN u1_slt4_reg_b14_b (.CK(bit_clk_pad_i), .D(n_10958), .Q(in_slt_432), .SO(in_slt_432), .SE(scan_enable), .SI(in_slt_410));
SDFFNSRN u1_slt6_reg_b14_b (.CK(bit_clk_pad_i), .D(n_10957), .Q(in_slt_454), .SO(in_slt_454), .SE(scan_enable), .SI(in_slt_432));
SDFFNSRN u1_slt2_reg_b14_b (.CK(bit_clk_pad_i), .D(n_10964), .Q(in_slt_840), .SO(in_slt_840), .SE(scan_enable), .SI(in_slt_454));
SDFFNSRN u1_sr_reg_b16_b (.CK(bit_clk_pad_i), .D(u1_sr_131), .Q(u1_sr_132), .SO(u1_sr_132), .SE(scan_enable), .SI(in_slt_840));
SDFFNSRN u1_slt2_reg_b13_b (.CK(bit_clk_pad_i), .D(n_10804), .Q(in_slt_839), .SO(in_slt_839), .SE(scan_enable), .SI(u1_sr_132));
SDFFNSRN u1_slt4_reg_b13_b (.CK(bit_clk_pad_i), .D(n_10802), .Q(in_slt_431), .SO(in_slt_431), .SE(scan_enable), .SI(in_slt_839));
SDFFNSRN u1_slt6_reg_b13_b (.CK(bit_clk_pad_i), .D(n_10800), .Q(in_slt_453), .SO(in_slt_453), .SE(scan_enable), .SI(in_slt_431));
SDFFNSRN u1_slt3_reg_b13_b (.CK(bit_clk_pad_i), .D(n_10803), .Q(in_slt_409), .SO(in_slt_409), .SE(scan_enable), .SI(in_slt_453));
SDFFNSRN u1_sr_reg_b15_b (.CK(bit_clk_pad_i), .D(u1_sr_130), .Q(u1_sr_131), .SO(u1_sr_131), .SE(scan_enable), .SI(in_slt_409));
SDFFNSRN u0_slt9_r_reg_b3_b (.CK(bit_clk_pad_i), .D(n_9953), .Q(u0_slt9_r_170), .SO(u0_slt9_r_170), .SE(scan_enable), .SI(u1_sr_131));
SDFFNSRN u1_slt6_reg_b12_b (.CK(bit_clk_pad_i), .D(n_9954), .Q(in_slt_452), .SO(in_slt_452), .SE(scan_enable), .SI(u0_slt9_r_170));
SDFFNSRN u1_slt0_reg_b12_b (.CK(bit_clk_pad_i), .D(n_9958), .Q(in_slt_739), .SO(in_slt_739), .SE(scan_enable), .SI(in_slt_452));
SDFFNSRN u1_slt2_reg_b12_b (.CK(bit_clk_pad_i), .D(n_9957), .Q(in_slt_838), .SO(in_slt_838), .SE(scan_enable), .SI(in_slt_739));
SDFFNSRN u1_slt3_reg_b12_b (.CK(bit_clk_pad_i), .D(n_9956), .Q(in_slt_408), .SO(in_slt_408), .SE(scan_enable), .SI(in_slt_838));
SDFFNSRN u1_slt4_reg_b12_b (.CK(bit_clk_pad_i), .D(n_9955), .Q(in_slt_430), .SO(in_slt_430), .SE(scan_enable), .SI(in_slt_408));
SDFFNSRN u1_sr_reg_b14_b (.CK(bit_clk_pad_i), .D(u1_sr_129), .Q(u1_sr_130), .SO(u1_sr_130), .SE(scan_enable), .SI(in_slt_430));
SDFFNSRN u1_slt4_reg_b11_b (.CK(bit_clk_pad_i), .D(n_9761), .Q(in_slt_429), .SO(in_slt_429), .SE(scan_enable), .SI(u1_sr_130));
SDFFNSRN u1_slt0_reg_b11_b (.CK(bit_clk_pad_i), .D(n_9765), .Q(in_slt_738), .SO(in_slt_738), .SE(scan_enable), .SI(in_slt_429));
SDFFNSRN u1_slt1_reg_b11_b (.CK(bit_clk_pad_i), .D(n_9764), .Q(in_slt_753), .SO(in_slt_753), .SE(scan_enable), .SI(in_slt_738));
SDFFNSRN u1_slt2_reg_b11_b (.CK(bit_clk_pad_i), .D(n_9763), .Q(in_slt_837), .SO(in_slt_837), .SE(scan_enable), .SI(in_slt_753));
SDFFNSRN u1_slt3_reg_b11_b (.CK(bit_clk_pad_i), .D(n_9762), .Q(in_slt_407), .SO(in_slt_407), .SE(scan_enable), .SI(in_slt_837));
SDFFNSRN u1_slt6_reg_b11_b (.CK(bit_clk_pad_i), .D(n_9760), .Q(in_slt_451), .SO(in_slt_451), .SE(scan_enable), .SI(in_slt_407));
SDFFNSRN u1_sr_reg_b13_b (.CK(bit_clk_pad_i), .D(u1_sr_128), .Q(u1_sr_129), .SO(u1_sr_129), .SE(scan_enable), .SI(in_slt_451));
SDFFNSRN u1_slt6_reg_b10_b (.CK(bit_clk_pad_i), .D(n_9618), .Q(in_slt_450), .SO(in_slt_450), .SE(scan_enable), .SI(u1_sr_129));
SDFFNSRN u1_slt2_reg_b10_b (.CK(bit_clk_pad_i), .D(n_9628), .Q(in_slt_836), .SO(in_slt_836), .SE(scan_enable), .SI(in_slt_450));
SDFFNSRN u1_slt1_reg_b10_b (.CK(bit_clk_pad_i), .D(n_9630), .Q(in_slt_752), .SO(in_slt_752), .SE(scan_enable), .SI(in_slt_836));
SDFFNSRN u1_slt4_reg_b10_b (.CK(bit_clk_pad_i), .D(n_9619), .Q(in_slt_428), .SO(in_slt_428), .SE(scan_enable), .SI(in_slt_752));
SDFFNSRN u1_slt3_reg_b10_b (.CK(bit_clk_pad_i), .D(n_9625), .Q(in_slt_406), .SO(in_slt_406), .SE(scan_enable), .SI(in_slt_428));
SDFFNSRN u0_slt9_r_reg_b2_b (.CK(bit_clk_pad_i), .D(n_9603), .Q(u0_slt9_r_169), .SO(u0_slt9_r_169), .SE(scan_enable), .SI(in_slt_406));
SDFFNSRN u1_sr_reg_b12_b (.CK(bit_clk_pad_i), .D(u1_sr_127), .Q(u1_sr_128), .SO(u1_sr_128), .SE(scan_enable), .SI(u0_slt9_r_169));
SDFFNSRN u1_slt2_reg_b9_b (.CK(bit_clk_pad_i), .D(n_9530), .Q(in_slt_835), .SO(in_slt_835), .SE(scan_enable), .SI(u1_sr_128));
SDFFNSRN u1_slt0_reg_b9_b (.CK(bit_clk_pad_i), .D(n_9531), .Q(in_slt_736), .SO(in_slt_736), .SE(scan_enable), .SI(in_slt_835));
SDFFNSRN u1_slt4_reg_b9_b (.CK(bit_clk_pad_i), .D(n_9528), .Q(in_slt_427), .SO(in_slt_427), .SE(scan_enable), .SI(in_slt_736));
SDFFNSRN u1_slt3_reg_b9_b (.CK(bit_clk_pad_i), .D(n_9529), .Q(in_slt_405), .SO(in_slt_405), .SE(scan_enable), .SI(in_slt_427));
SDFFNSRN u1_slt6_reg_b9_b (.CK(bit_clk_pad_i), .D(n_9527), .Q(in_slt_449), .SO(in_slt_449), .SE(scan_enable), .SI(in_slt_405));
SDFFNSRN u1_sr_reg_b11_b (.CK(bit_clk_pad_i), .D(u1_sr_126), .Q(u1_sr_127), .SO(u1_sr_127), .SE(scan_enable), .SI(in_slt_449));
SDFFNSRN u1_slt6_reg_b8_b (.CK(bit_clk_pad_i), .D(n_9353), .Q(in_slt_448), .SO(in_slt_448), .SE(scan_enable), .SI(u1_sr_127));
SDFFNSRN u1_slt2_reg_b8_b (.CK(bit_clk_pad_i), .D(n_9356), .Q(in_slt_834), .SO(in_slt_834), .SE(scan_enable), .SI(in_slt_448));
SDFFNSRN u1_slt1_reg_b8_b (.CK(bit_clk_pad_i), .D(n_9357), .Q(in_slt_750), .SO(in_slt_750), .SE(scan_enable), .SI(in_slt_834));
SDFFNSRN u1_slt4_reg_b8_b (.CK(bit_clk_pad_i), .D(n_9354), .Q(in_slt_426), .SO(in_slt_426), .SE(scan_enable), .SI(in_slt_750));
SDFFNSRN u1_slt3_reg_b8_b (.CK(bit_clk_pad_i), .D(n_9355), .Q(in_slt_404), .SO(in_slt_404), .SE(scan_enable), .SI(in_slt_426));
SDFFNSRN u1_sr_reg_b10_b (.CK(bit_clk_pad_i), .D(u1_sr_125), .Q(u1_sr_126), .SO(u1_sr_126), .SE(scan_enable), .SI(in_slt_404));
SDFFNSRN u1_slt1_reg_b7_b (.CK(bit_clk_pad_i), .D(n_8258), .Q(in_slt_749), .SO(in_slt_749), .SE(scan_enable), .SI(u1_sr_126));
SDFFNSRN u1_slt2_reg_b7_b (.CK(bit_clk_pad_i), .D(n_8257), .Q(in_slt_833), .SO(in_slt_833), .SE(scan_enable), .SI(in_slt_749));
SDFFNSRN u1_slt4_reg_b7_b (.CK(bit_clk_pad_i), .D(n_8255), .Q(in_slt_425), .SO(in_slt_425), .SE(scan_enable), .SI(in_slt_833));
SDFFNSRN u1_slt3_reg_b7_b (.CK(bit_clk_pad_i), .D(n_8256), .Q(in_slt_403), .SO(in_slt_403), .SE(scan_enable), .SI(in_slt_425));
SDFFNSRN u0_slt9_r_reg_b1_b (.CK(bit_clk_pad_i), .D(n_8211), .Q(u0_slt9_r_168), .SO(u0_slt9_r_168), .SE(scan_enable), .SI(in_slt_403));
SDFFNSRN u1_slt6_reg_b7_b (.CK(bit_clk_pad_i), .D(n_8254), .Q(in_slt_447), .SO(in_slt_447), .SE(scan_enable), .SI(u0_slt9_r_168));
SDFFNSRN u1_sr_reg_b9_b (.CK(bit_clk_pad_i), .D(u1_sr_124), .Q(u1_sr_125), .SO(u1_sr_125), .SE(scan_enable), .SI(in_slt_447));
SDFFNSRN u1_slt3_reg_b6_b (.CK(bit_clk_pad_i), .D(n_7509), .Q(in_slt_402), .SO(in_slt_402), .SE(scan_enable), .SI(u1_sr_125));
SDFFNSRN u1_slt1_reg_b6_b (.CK(bit_clk_pad_i), .D(n_7507), .Q(in_slt_748), .SO(in_slt_748), .SE(scan_enable), .SI(in_slt_402));
SDFFNSRN u1_slt2_reg_b6_b (.CK(bit_clk_pad_i), .D(n_7510), .Q(in_slt_832), .SO(in_slt_832), .SE(scan_enable), .SI(in_slt_748));
SDFFNSRN u1_slt4_reg_b6_b (.CK(bit_clk_pad_i), .D(n_7511), .Q(in_slt_424), .SO(in_slt_424), .SE(scan_enable), .SI(in_slt_832));
SDFFNSRN u1_slt6_reg_b6_b (.CK(bit_clk_pad_i), .D(n_7508), .Q(in_slt_446), .SO(in_slt_446), .SE(scan_enable), .SI(in_slt_424));
SDFFNSRN u1_sr_reg_b8_b (.CK(bit_clk_pad_i), .D(u1_sr_123), .Q(u1_sr_124), .SO(u1_sr_124), .SE(scan_enable), .SI(in_slt_446));
SDFFNSRN u1_slt1_reg_b5_b (.CK(bit_clk_pad_i), .D(n_7359), .Q(in_slt_747), .SO(in_slt_747), .SE(scan_enable), .SI(u1_sr_124));
SDFFNSRN u1_slt2_reg_b5_b (.CK(bit_clk_pad_i), .D(n_7360), .Q(in_slt_831), .SO(in_slt_831), .SE(scan_enable), .SI(in_slt_747));
SDFFNSRN u1_slt4_reg_b5_b (.CK(bit_clk_pad_i), .D(n_7362), .Q(in_slt_423), .SO(in_slt_423), .SE(scan_enable), .SI(in_slt_831));
SDFFNSRN u1_slt3_reg_b5_b (.CK(bit_clk_pad_i), .D(n_7358), .Q(in_slt_401), .SO(in_slt_401), .SE(scan_enable), .SI(in_slt_423));
SDFFNSRN u1_slt6_reg_b5_b (.CK(bit_clk_pad_i), .D(n_7361), .Q(in_slt_445), .SO(in_slt_445), .SE(scan_enable), .SI(in_slt_401));
SDFFNSRN u1_sr_reg_b7_b (.CK(bit_clk_pad_i), .D(u1_sr_122), .Q(u1_sr_123), .SO(u1_sr_123), .SE(scan_enable), .SI(in_slt_445));
SDFFNSRN u0_slt9_r_reg_b0_b (.CK(bit_clk_pad_i), .D(n_7231), .Q(u0_slt9_r), .SO(u0_slt9_r), .SE(scan_enable), .SI(u1_sr_123));
SDFFNSRN u1_slt2_reg_b4_b (.CK(bit_clk_pad_i), .D(n_7144), .Q(in_slt_830), .SO(in_slt_830), .SE(scan_enable), .SI(u0_slt9_r));
SDFFNSRN u1_slt3_reg_b4_b (.CK(bit_clk_pad_i), .D(n_7156), .Q(in_slt_400), .SO(in_slt_400), .SE(scan_enable), .SI(in_slt_830));
SDFFNSRN u1_slt4_reg_b4_b (.CK(bit_clk_pad_i), .D(n_7155), .Q(in_slt_422), .SO(in_slt_422), .SE(scan_enable), .SI(in_slt_400));
SDFFNSRN u1_slt6_reg_b4_b (.CK(bit_clk_pad_i), .D(n_7154), .Q(in_slt_444), .SO(in_slt_444), .SE(scan_enable), .SI(in_slt_422));
SDFFNSRN u1_sr_reg_b6_b (.CK(bit_clk_pad_i), .D(u1_sr_121), .Q(u1_sr_122), .SO(u1_sr_122), .SE(scan_enable), .SI(in_slt_444));
SDFFNSRN u1_slt3_reg_b0_b (.CK(bit_clk_pad_i), .D(n_6731), .Q(in_slt3), .SO(in_slt3), .SE(scan_enable), .SI(u1_sr_122));
SDFFN u2_cnt_reg_b7_b (.CK(bit_clk_pad_i), .D(n_6066), .Q(n_1212), .SO(n_1212), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(in_slt3));
SDFFNSRN u1_slt3_reg_b2_b (.CK(bit_clk_pad_i), .D(n_6730), .Q(in_slt_398), .SO(in_slt_398), .SE(scan_enable), .SI(n_1212));
SDFFNSRN u1_slt3_reg_b1_b (.CK(bit_clk_pad_i), .D(n_6732), .Q(in_slt_397), .SO(in_slt_397), .SE(scan_enable), .SI(in_slt_398));
SDFFNSRN u1_slt4_reg_b1_b (.CK(bit_clk_pad_i), .D(n_6727), .Q(in_slt_419), .SO(in_slt_419), .SE(scan_enable), .SI(in_slt_397));
SDFFNSRN u1_slt6_reg_b1_b (.CK(bit_clk_pad_i), .D(n_6723), .Q(in_slt_441), .SO(in_slt_441), .SE(scan_enable), .SI(in_slt_419));
SDFFNSRN u1_slt6_reg_b2_b (.CK(bit_clk_pad_i), .D(n_6722), .Q(in_slt_442), .SO(in_slt_442), .SE(scan_enable), .SI(in_slt_441));
SDFFNSRN u1_slt6_reg_b3_b (.CK(bit_clk_pad_i), .D(n_6721), .Q(in_slt_443), .SO(in_slt_443), .SE(scan_enable), .SI(in_slt_442));
SDFFNSRN u1_slt6_reg_b0_b (.CK(bit_clk_pad_i), .D(n_6724), .Q(in_slt6), .SO(in_slt6), .SE(scan_enable), .SI(in_slt_443));
SDFFNSRN u1_slt4_reg_b3_b (.CK(bit_clk_pad_i), .D(n_6725), .Q(in_slt_421), .SO(in_slt_421), .SE(scan_enable), .SI(in_slt6));
SDFFNSRN u1_slt3_reg_b3_b (.CK(bit_clk_pad_i), .D(n_6729), .Q(in_slt_399), .SO(in_slt_399), .SE(scan_enable), .SI(in_slt_421));
SDFFNSRN u1_slt4_reg_b2_b (.CK(bit_clk_pad_i), .D(n_6726), .Q(in_slt_420), .SO(in_slt_420), .SE(scan_enable), .SI(in_slt_399));
SDFFNSRN u1_slt4_reg_b0_b (.CK(bit_clk_pad_i), .D(n_6728), .Q(in_slt4), .SO(in_slt4), .SE(scan_enable), .SI(in_slt_420));
SDFFN u2_cnt_reg_b1_b (.CK(bit_clk_pad_i), .D(n_5821), .Q(n_866), .SO(n_866), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(in_slt4));
SDFFNSRN u1_sr_reg_b5_b (.CK(bit_clk_pad_i), .D(u1_sr_120), .Q(u1_sr_121), .SO(u1_sr_121), .SE(scan_enable), .SI(n_866));
SDFFN u2_cnt_reg_b4_b (.CK(bit_clk_pad_i), .D(n_6058), .Q(u2_cnt_b4_b), .SO(u2_cnt_b4_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u1_sr_121));
SDFFN u2_cnt_reg_b3_b (.CK(bit_clk_pad_i), .D(n_6052), .Q(u2_cnt_b3_b), .SO(u2_cnt_b3_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u2_cnt_b4_b));
SDFFN u2_cnt_reg_b5_b (.CK(bit_clk_pad_i), .D(n_5741), .Q(u2_cnt_b5_b), .SO(u2_cnt_b5_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u2_cnt_b3_b));
SDFFN u2_cnt_reg_b6_b (.CK(bit_clk_pad_i), .D(n_5889), .Q(u2_cnt_b6_b), .SO(u2_cnt_b6_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u2_cnt_b5_b));
SDFFN u2_cnt_reg_b0_b (.CK(bit_clk_pad_i), .D(n_5822), .Q(n_1773), .SO(n_1773), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u2_cnt_b6_b));
SDFFN u2_cnt_reg_b2_b (.CK(bit_clk_pad_i), .D(n_5820), .Q(u2_cnt_b2_b), .SO(u2_cnt_b2_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(n_1773));
SDFFNSRN u2_valid_reg (.CK(bit_clk_pad_i), .D(n_5611), .Q(valid), .SO(valid), .SE(scan_enable), .SI(u2_cnt_b2_b));
SDFFNSRN u2_in_valid_reg_b0_b (.CK(bit_clk_pad_i), .D(n_5593), .Q(in_valid), .SO(in_valid), .SE(scan_enable), .SI(valid));
SDFFNSRN u1_sr_reg_b4_b (.CK(bit_clk_pad_i), .D(u1_sr_119), .Q(u1_sr_120), .SO(u1_sr_120), .SE(scan_enable), .SI(in_valid));
SDFFNSRN u2_in_valid_reg_b2_b (.CK(bit_clk_pad_i), .D(n_5432), .Q(in_valid_9), .SO(in_valid_9), .SE(scan_enable), .SI(u1_sr_120));
SDFFNSRN u2_sync_beat_reg (.CK(bit_clk_pad_i), .D(n_5441), .Q(u2_sync_beat), .SO(u2_sync_beat), .SE(scan_enable), .SI(in_valid_9));
SDFFNSRN u2_ld_reg (.CK(bit_clk_pad_i), .D(n_4833), .Q(n_6734), .SO(n_6734), .SE(scan_enable), .SI(u2_sync_beat));
SDFFNSRN u2_out_le_reg_b1_b (.CK(bit_clk_pad_i), .D(n_4831), .Q(out_le_180), .SO(out_le_180), .SE(scan_enable), .SI(n_6734));
SDFFNSRN u2_in_valid_reg_b1_b (.CK(bit_clk_pad_i), .D(n_4840), .Q(in_valid_8), .SO(in_valid_8), .SE(scan_enable), .SI(out_le_180));
SDFFN u2_out_le_reg_b2_b (.CK(bit_clk_pad_i), .D(n_4077), .Q(out_le_181), .SO(out_le_181), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(in_valid_8));
SDFFN u2_out_le_reg_b4_b (.CK(bit_clk_pad_i), .D(n_4096), .Q(out_le_183), .SO(out_le_183), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(out_le_181));
SDFFN u2_out_le_reg_b5_b (.CK(bit_clk_pad_i), .D(n_4095), .Q(out_le_184), .SO(out_le_184), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(out_le_183));
SDFFN u2_out_le_reg_b3_b (.CK(bit_clk_pad_i), .D(n_4107), .Q(out_le_182), .SO(out_le_182), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(out_le_184));
SDFFNSRN u2_out_le_reg_b0_b (.CK(bit_clk_pad_i), .D(n_3984), .Q(out_le), .SO(out_le), .SE(scan_enable), .SI(out_le_182));
SDFFNSRN u1_sr_reg_b3_b (.CK(bit_clk_pad_i), .D(u1_sr_118), .Q(u1_sr_119), .SO(u1_sr_119), .SE(scan_enable), .SI(out_le));
SDFFNSRN u1_sr_reg_b2_b (.CK(bit_clk_pad_i), .D(u1_sr_117), .Q(u1_sr_118), .SO(u1_sr_118), .SE(scan_enable), .SI(u1_sr_119));
SDFFNSRN u1_sr_reg_b1_b (.CK(bit_clk_pad_i), .D(u1_sr), .Q(u1_sr_117), .SO(u1_sr_117), .SE(scan_enable), .SI(u1_sr_118));
SDFFNSRN u1_sr_reg_b0_b (.CK(bit_clk_pad_i), .D(u1_sdata_in_r), .Q(u1_sr), .SO(u1_sr), .SE(scan_enable), .SI(u1_sr_117));
// scan chain ends here

 buf1 BUFbread(scan_data_out, u1_sr);
MX2X1 g29860(.A (n_208), .B (u0_slt9_r_182), .S0 (n_11395), .Y(n_11214));
MX2X1 g29862(.A (n_297), .B (u0_slt9_r_181), .S0 (n_11319), .Y(n_11213));
MX2X1 g29688(.A (n_10790), .B (u0_slt4_r_73), .S0 (n_6710), .Y(n_11312));
MX2X1 g29866(.A (n_203), .B (u0_slt9_r_179), .S0 (n_11389), .Y(n_11211));
MX2X1 g29684(.A (n_373), .B (u0_slt4_r_75), .S0 (n_11319), .Y(n_11314));
MX2X1 g29686(.A (n_10788), .B (u0_slt4_r_74), .S0 (n_11389), .Y(n_11313));
MX2X1 g29680(.A (n_370), .B (u0_slt4_r_77), .S0 (n_11389), .Y(n_11317));
MX2X1 g29682(.A (n_380), .B (u0_slt4_r_76), .S0 (n_7042), .Y(n_11315));
INVX1 g41880(.A (u2_cnt_b3_b ), .Y (n_698));
MX2X1 g29864(.A (n_263), .B (u0_slt9_r_180), .S0 (n_11389), .Y(n_11212));
MX2X1 g29868(.A (n_152), .B (u0_slt9_r_178), .S0 (n_7042), .Y(n_11210));
AOI21X1 g40392(.A0 (n_688), .A1 (n_866), .B0 (n_1824), .Y (n_1928));
AOI21X1 g36614(.A0 (n_2572), .A1 (u2_cnt_b6_b ), .B0 (n_1212), .Y(n_5430));
INVX1 g42138(.A (out_slt3), .Y (n_251));
MX2X1 g29808(.A (n_10990), .B (u0_slt7_r_130), .S0 (n_11395), .Y(n_11243));
MX2X1 g29802(.A (n_201), .B (u0_slt7_r_133), .S0 (n_6710), .Y(n_11246));
MX2X1 g29800(.A (n_217), .B (u0_slt7_r_134), .S0 (n_11319), .Y(n_11247));
MX2X1 g29806(.A (n_10988), .B (u0_slt7_r_131), .S0 (n_11389), .Y(n_11244));
MX2X1 g29804(.A (n_335), .B (u0_slt7_r_132), .S0 (n_11389), .Y(n_11245));
INVX1 g42875(.A (out_slt_67), .Y (n_10976));
INVX1 g42724(.A (out_slt_146), .Y (n_352));
INVX1 g42723(.A (out_slt_102), .Y (n_361));
NAND2X1 g35839(.A (n_4826), .B (n_6057), .Y (n_5741));
NOR2X1 g35855(.A (n_1823), .B (n_1469), .Y (n_4107));
OR2X1 g35676(.A (n_1087), .B (n_7042), .Y (n_7043));
INVX1 g42446(.A (out_slt_175), .Y (n_208));
INVX1 g42114(.A (out_slt_168), .Y (n_183));
MX2X1 g29824(.A (n_228), .B (u0_slt8_r_161), .S0 (n_11319), .Y(n_11235));
MX2X1 g29826(.A (n_76), .B (u0_slt8_r_160), .S0 (n_6710), .Y(n_11234));
MX2X1 g29820(.A (n_79), .B (u0_slt8_r_163), .S0 (n_11319), .Y(n_11237));
MX2X1 g29822(.A (n_237), .B (u0_slt8_r_162), .S0 (n_11395), .Y(n_11236));
MX2X1 g29828(.A (n_212), .B (u0_slt8_r_159), .S0 (n_11319), .Y(n_11233));
MX2X1 g30130(.A (in_slt_739), .B (u1_sr_128), .S0 (out_le), .Y(n_9958));
MX2X1 g29536(.A (crac_out_867), .B (u0_slt1_r_32), .S0 (n_11389), .Y(n_11416));
MX2X1 g29534(.A (crac_out_876), .B (u0_slt1_r_33), .S0 (n_11389), .Y(n_11417));
AND2X1 g29532(.A (u0_slt1_r_34), .B (n_11395), .Y (n_11418));
AND2X1 g29530(.A (u0_slt0_r), .B (n_11395), .Y (n_11419));
MX2X1 g29538(.A (crac_out_866), .B (u0_slt1_r_31), .S0 (n_11319), .Y(n_11414));
MX2X1 g29778(.A (n_163), .B (u0_slt7_r_145), .S0 (n_11319), .Y(n_11258));
MX2X1 g29774(.A (n_299), .B (u0_slt7_r_147), .S0 (n_11389), .Y(n_11262));
INVX1 g41790(.A (out_slt_145), .Y (n_280));
INVX4 g35762(.A (n_7038), .Y (n_11395));
BUFX3 g35760(.A (n_6734), .Y (n_6710));
INVX1 g41794(.A (crac_out_848), .Y (n_71));
INVX1 g35769(.A (n_7042), .Y (n_7038));
AND2X1 g29708(.A (u0_slt5_r_102), .B (n_11395), .Y (n_11301));
AND2X1 g29704(.A (u0_slt5_r_104), .B (n_11395), .Y (n_11303));
AND2X1 g29706(.A (u0_slt5_r_103), .B (n_11395), .Y (n_11302));
AND2X1 g29700(.A (u0_slt5_r_106), .B (n_11395), .Y (n_11305));
AND2X1 g29702(.A (u0_slt5_r_105), .B (n_11395), .Y (n_11304));
OR2X1 g36306(.A (n_2597), .B (n_1212), .Y (n_4840));
MX2X1 g31309(.A (u1_sr_126), .B (in_slt_428), .S0 (out_le_183), .Y(n_9619));
MX2X1 g31300(.A (u1_sr_126), .B (in_slt_406), .S0 (out_le_182), .Y(n_9625));
INVX1 g41978(.A (out_slt_162), .Y (n_9952));
INVX1 g42686(.A (out_slt_129), .Y (n_265));
INVX1 g42468(.A (crac_out_858), .Y (n_179));
MX2X1 g35379(.A (u1_sr_119), .B (in_slt_443), .S0 (out_le_184), .Y(n_6721));
MX2X1 g35378(.A (u1_sr_118), .B (in_slt_442), .S0 (out_le_184), .Y(n_6722));
MX2X1 g35371(.A (u1_sr), .B (in_slt4), .S0 (out_le_183), .Y (n_6728));
MX2X1 g35370(.A (u1_sr_121), .B (in_slt_401), .S0 (out_le_182), .Y(n_7358));
MX2X1 g35373(.A (u1_sr_118), .B (in_slt_420), .S0 (out_le_183), .Y(n_6726));
MX2X1 g35372(.A (u1_sr_117), .B (in_slt_419), .S0 (out_le_183), .Y(n_6727));
MX2X1 g35375(.A (u1_sr_120), .B (in_slt_422), .S0 (out_le_183), .Y(n_7155));
MX2X1 g35377(.A (u1_sr_117), .B (in_slt_441), .S0 (out_le_184), .Y(n_6723));
NAND3X1 g36565(.A (n_1822), .B (n_1824), .C (n_684), .Y (n_1825));
AND2X1 g29511(.A (u0_slt0_r_9), .B (n_7042), .Y (n_11431));
MX2X1 g29513(.A (out_slt_20), .B (u0_slt0_r_8), .S0 (n_11319), .Y(n_11430));
MX2X1 g29515(.A (out_slt_19), .B (u0_slt0_r_7), .S0 (n_11389), .Y(n_11429));
MX2X1 g29517(.A (out_slt_18), .B (u0_slt0_r_6), .S0 (n_11389), .Y(n_11428));
AOI21X1 g36449(.A0 (n_3965), .A1 (n_3995), .B0 (n_4079), .Y (n_5611));
INVX1 g42096(.A (out_slt_80), .Y (n_281));
INVX1 g42094(.A (out_slt_164), .Y (n_359));
MX2X1 g29876(.A (n_160), .B (u0_slt9_r_174), .S0 (n_11389), .Y(n_11205));
MX2X1 g29874(.A (n_183), .B (u0_slt9_r_175), .S0 (n_11389), .Y(n_11206));
AND2X1 g29696(.A (u0_slt5_r_108), .B (n_11395), .Y (n_11307));
AND2X1 g29694(.A (u0_slt5_r_109), .B (n_11395), .Y (n_11308));
INVX1 g36613(.A (n_5430), .Y (n_5593));
INVX8 g35740(.A (n_6999), .Y (n_11389));
INVX2 g35744(.A (n_6710), .Y (n_6999));
AND2X1 g29726(.A (u0_slt5_r_93), .B (n_11395), .Y (n_11292));
AND2X1 g29724(.A (u0_slt5_r_94), .B (n_11395), .Y (n_11293));
AND2X1 g29722(.A (u0_slt5_r_95), .B (n_11395), .Y (n_11294));
AND2X1 g29720(.A (u0_slt5_r_96), .B (n_11395), .Y (n_11295));
AND2X1 g29728(.A (u0_slt5_r_92), .B (n_11395), .Y (n_11291));
INVX1 g42666(.A (crac_out_846), .Y (n_227));
INVX1 g42661(.A (out_slt_158), .Y (n_86));
NAND2X1 g35843(.A (n_3996), .B (n_4832), .Y (n_5441));
INVX1 g42401(.A (n_1212), .Y (n_456));
INVX1 g42407(.A (u2_cnt_b5_b ), .Y (n_701));
NAND2X1 g35840(.A (n_4825), .B (n_6057), .Y (n_5889));
MX2X1 g29578(.A (n_179), .B (u0_slt2_r_50), .S0 (n_11389), .Y(n_11387));
AND2X1 g29572(.A (u0_slt2_r_53), .B (n_11395), .Y (n_11391));
AND2X1 g29570(.A (u0_slt1_r), .B (n_11395), .Y (n_11392));
MX2X1 g29576(.A (n_177), .B (u0_slt2_r_51), .S0 (n_11319), .Y(n_11388));
MX2X1 g29574(.A (n_170), .B (u0_slt2_r_52), .S0 (n_11389), .Y(n_11390));
INVX1 g42340(.A (out_slt_77), .Y (n_195));
INVX1 g35720(.A (n_2631), .Y (n_2632));
MX2X1 g29740(.A (n_113), .B (u0_slt6_r_125), .S0 (n_11319), .Y(n_11284));
MX2X1 g29742(.A (n_101), .B (u0_slt6_r_124), .S0 (n_11389), .Y(n_11283));
MX2X1 g29961(.A (u1_sr_132), .B (in_slt_456), .S0 (out_le_184), .Y(n_11166));
MX2X1 g29744(.A (n_261), .B (u0_slt6_r_123), .S0 (n_7042), .Y(n_11281));
MX2X1 g29746(.A (n_300), .B (u0_slt6_r_122), .S0 (n_11319), .Y(n_11280));
MX2X1 g29748(.A (n_84), .B (u0_slt6_r_121), .S0 (n_11319), .Y(n_11279));
NAND2X1 g37471(.A (n_1784), .B (u2_cnt_b5_b ), .Y (n_1785));
NAND2X1 g37472(.A (n_2592), .B (n_688), .Y (n_1782));
OR2X1 g37473(.A (n_3964), .B (n_2596), .Y (n_3965));
MX2X1 g29898(.A (u1_sr_135), .B (in_slt_437), .S0 (out_le_183), .Y(n_11200));
XOR2X1 g34903(.A (n_1212), .B (n_4103), .Y (n_5635));
MX2X1 g29880(.A (n_372), .B (u0_slt9_r_172), .S0 (n_6710), .Y(n_11203));
AND2X1 g29554(.A (u0_slt1_r_23), .B (n_11395), .Y (n_11403));
AND2X1 g29556(.A (u0_slt1_r_22), .B (n_7042), .Y (n_11401));
AND2X1 g29550(.A (u0_slt1_r_25), .B (n_11395), .Y (n_11406));
AND2X1 g29552(.A (u0_slt1_r_24), .B (n_11395), .Y (n_11404));
AND2X1 g29558(.A (u0_slt1_r_21), .B (n_11395), .Y (n_11400));
NAND3X1 g39333(.A (n_698), .B (u2_cnt_b5_b ), .C (n_456), .Y (n_1486));
INVX1 g42364(.A (out_slt_18), .Y (n_1100));
INVX1 g43016(.A (out_slt_143), .Y (n_10981));
INVX1 g43012(.A (out_slt_166), .Y (n_191));
MX2X1 g34070(.A (u1_sr_123), .B (in_slt_749), .S0 (out_le_180), .Y(n_8258));
MX2X1 g29768(.A (n_10785), .B (u0_slt6_r_111), .S0 (n_11319), .Y(n_11266));
MX2X1 g29762(.A (n_262), .B (u0_slt6_r_114), .S0 (n_11319), .Y(n_11269));
MX2X1 g29760(.A (n_234), .B (u0_slt6_r_115), .S0 (n_11319), .Y(n_11270));
MX2X1 g29766(.A (n_10783), .B (u0_slt6_r_112), .S0 (n_11389), .Y(n_11267));
MX2X1 g29764(.A (n_304), .B (u0_slt6_r_113), .S0 (n_11389), .Y(n_11268));
INVX1 g42193(.A (crac_out_850), .Y (n_311));
MX2X1 g34914(.A (u1_sr_122), .B (in_slt_446), .S0 (out_le_184), .Y(n_7508));
MX2X1 g34915(.A (u1_sr_122), .B (in_slt_748), .S0 (out_le_180), .Y(n_7507));
AND2X1 g41536(.A (n_701), .B (n_2596), .Y (n_2571));
INVX1 g41859(.A (out_slt_73), .Y (n_341));
INVX1 g42818(.A (u2_cnt_b2_b ), .Y (n_684));
INVX1 g42819(.A (out_slt_81), .Y (n_109));
INVX1 g42971(.A (crac_out_856), .Y (n_138));
INVX1 g41779(.A (out_slt_66), .Y (n_10978));
INVX1 g42924(.A (out_slt_173), .Y (n_263));
AOI21X1 g36741(.A0 (n_2602), .A1 (u2_cnt_b6_b ), .B0 (n_2603), .Y(n_4825));
MX2X1 g30034(.A (u1_sr_130), .B (in_slt_454), .S0 (out_le_184), .Y(n_10957));
MX2X1 g30031(.A (u1_sr_130), .B (in_slt_840), .S0 (out_le_181), .Y(n_10964));
MX2X1 g30033(.A (u1_sr_130), .B (in_slt_432), .S0 (out_le_183), .Y(n_10958));
MX2X1 g30032(.A (u1_sr_130), .B (in_slt_410), .S0 (out_le_182), .Y(n_10961));
MX2X1 g29598(.A (n_71), .B (u0_slt2_r_40), .S0 (n_11319), .Y(n_11373));
MX2X1 g29590(.A (n_357), .B (u0_slt2_r_44), .S0 (n_11395), .Y(n_11378));
MX2X1 g29592(.A (n_149), .B (u0_slt2_r_43), .S0 (n_11389), .Y(n_11377));
MX2X1 g29594(.A (n_311), .B (u0_slt2_r_42), .S0 (n_11319), .Y(n_11376));
MX2X1 g29596(.A (n_130), .B (u0_slt2_r_41), .S0 (n_11319), .Y(n_11375));
MX2X1 g29616(.A (n_16), .B (u0_slt3_r_70), .S0 (n_11389), .Y(n_11361));
MX2X1 g34912(.A (u1_sr_122), .B (in_slt_832), .S0 (out_le_181), .Y(n_7510));
MX2X1 g34913(.A (u1_sr_122), .B (in_slt_402), .S0 (out_le_182), .Y(n_7509));
INVX1 g42018(.A (out_slt_78), .Y (n_267));
NOR2X1 g35835(.A (n_1825), .B (n_1486), .Y (n_4096));
INVX1 g43054(.A (out_slt6), .Y (n_223));
INVX1 g41930(.A (out_slt_136), .Y (n_134));
MX2X1 g29674(.A (n_394), .B (u0_slt4_r_80), .S0 (n_11319), .Y(n_11321));
MX2X1 g29676(.A (n_391), .B (u0_slt4_r_79), .S0 (n_11319), .Y(n_11320));
MX2X1 g29670(.A (n_321), .B (u0_slt4_r_82), .S0 (n_11389), .Y(n_11324));
MX2X1 g29672(.A (n_320), .B (u0_slt4_r_81), .S0 (n_6710), .Y(n_11323));
MX2X1 g29678(.A (n_351), .B (u0_slt4_r_78), .S0 (n_7042), .Y(n_11318));
INVX1 g42831(.A (out_slt_123), .Y (n_10990));
INVX1 g42957(.A (out_slt_161), .Y (n_9602));
NOR2X1 g40883(.A (n_688), .B (n_866), .Y (n_1824));
INVX1 g42484(.A (out_slt_101), .Y (n_295));
INVX1 g42487(.A (out_slt_128), .Y (n_363));
INVX1 g42489(.A (out_slt_157), .Y (n_240));
INVX1 g42226(.A (crac_out_859), .Y (n_177));
INVX1 g42222(.A (out_slt_178), .Y (n_383));
INVX1 g42799(.A (out_slt_138), .Y (n_163));
NAND4X1 g37598(.A (n_1253), .B (n_1227), .C (u2_cnt_b4_b ), .D(u2_cnt_b5_b ), .Y (n_2602));
MX2X1 g31825(.A (n_9602), .B (u0_slt9_r_168), .S0 (n_11319), .Y(n_9603));
MX2X1 g31821(.A (u1_sr_125), .B (in_slt_835), .S0 (out_le_181), .Y(n_9530));
MX2X1 g31820(.A (in_slt_736), .B (u1_sr_125), .S0 (out_le), .Y(n_9531));
MX2X1 g31823(.A (u1_sr_125), .B (in_slt_427), .S0 (out_le_183), .Y(n_9528));
MX2X1 g31822(.A (u1_sr_125), .B (in_slt_405), .S0 (out_le_182), .Y(n_9529));
INVX1 g37371(.A (n_2593), .Y (n_3984));
INVX1 g42032(.A (out_slt_121), .Y (n_102));
INVX1 g42035(.A (out_slt_83), .Y (n_329));
INVX1 g43075(.A (u2_cnt_b6_b ), .Y (n_711));
MX2X1 g29658(.A (n_396), .B (u0_slt4_r_88), .S0 (n_6710), .Y(n_11332));
MX2X1 g29656(.A (n_295), .B (u0_slt4_r_89), .S0 (n_6710), .Y(n_11333));
MX2X1 g29654(.A (n_361), .B (u0_slt4_r_90), .S0 (n_11389), .Y(n_11334));
MX2X1 g29652(.A (n_251), .B (u0_slt4_r_91), .S0 (n_11319), .Y(n_11336));
MX2X1 g29650(.A (n_220), .B (u0_slt3_r), .S0 (n_11319), .Y (n_11338));
INVX1 g42857(.A (out_slt_169), .Y (n_308));
INVX1 g42854(.A (out_slt_156), .Y (n_79));
INVX1 g36561(.A (n_4832), .Y (n_4833));
AND2X1 g36560(.A (n_4000), .B (n_1212), .Y (n_5432));
NOR2X1 g36563(.A (n_1114), .B (n_2604), .Y (n_4831));
NAND4X1 g36562(.A (n_2378), .B (n_698), .C (n_2596), .D (n_4079), .Y(n_4832));
INVX1 g42933(.A (crac_out_857), .Y (n_338));
INVX1 g42209(.A (out_slt_110), .Y (n_266));
MX2X1 g30079(.A (u1_sr_129), .B (in_slt_409), .S0 (out_le_182), .Y(n_10803));
MX2X1 g30078(.A (u1_sr_129), .B (in_slt_839), .S0 (out_le_181), .Y(n_10804));
INVX1 g41865(.A (crac_out_860), .Y (n_170));
NAND2X1 g37578(.A (n_1520), .B (n_2571), .Y (n_2572));
AND2X1 g38955(.A (n_701), .B (n_3995), .Y (n_4079));
NAND3X1 g37594(.A (n_1519), .B (n_1773), .C (u2_cnt_b4_b ), .Y(n_1774));
INVX1 g35782(.A (n_6734), .Y (n_7003));
NOR2X1 g38951(.A (n_1114), .B (u2_cnt_b2_b ), .Y (n_2592));
INVX1 g43099(.A (out_slt_74), .Y (n_389));
INVX1 g43091(.A (out_slt_113), .Y (n_287));
INVX1 g41903(.A (out_slt_170), .Y (n_302));
MX2X1 g29638(.A (n_230), .B (u0_slt3_r_59), .S0 (n_11319), .Y(n_11347));
MX2X1 g29630(.A (n_398), .B (u0_slt3_r_63), .S0 (n_11395), .Y(n_11352));
MX2X1 g29632(.A (n_389), .B (u0_slt3_r_62), .S0 (n_11395), .Y(n_11351));
MX2X1 g29634(.A (n_341), .B (u0_slt3_r_61), .S0 (n_6710), .Y(n_11349));
MX2X1 g29636(.A (n_82), .B (u0_slt3_r_60), .S0 (n_11319), .Y(n_11348));
INVX1 g42793(.A (out_slt_122), .Y (n_22));
INVX1 g42267(.A (crac_out_849), .Y (n_130));
INVX1 g41974(.A (out_slt_72), .Y (n_82));
INVX1 g41977(.A (out_slt_115), .Y (n_300));
INVX1 g42075(.A (out_slt_65), .Y (n_220));
INVX1 g42070(.A (out_slt_159), .Y (n_328));
INVX1 g42072(.A (out_slt_108), .Y (n_234));
INVX1 g41837(.A (u2_cnt_b4_b ), .Y (n_2596));
INVX1 g41831(.A (out_slt_105), .Y (n_10783));
AND2X1 g29612(.A (u0_slt3_r_72), .B (n_11395), .Y (n_11364));
AND2X1 g29610(.A (u0_slt2_r), .B (n_7042), .Y (n_11365));
MX2X1 g29614(.A (n_329), .B (u0_slt3_r_71), .S0 (n_11389), .Y(n_11363));
MX2X1 g29618(.A (n_109), .B (u0_slt3_r_69), .S0 (n_11319), .Y(n_11360));
MX2X1 g31298(.A (u1_sr_126), .B (in_slt_836), .S0 (out_le_181), .Y(n_9628));
MX2X1 g31294(.A (u1_sr_126), .B (in_slt_752), .S0 (out_le_180), .Y(n_9630));
INVX1 g42119(.A (out_slt4), .Y (n_397));
INVX1 g42118(.A (out_slt_96), .Y (n_330));
INVX1 g41914(.A (out_slt_167), .Y (n_160));
NOR2X1 g40829(.A (u2_cnt_b4_b ), .B (n_711), .Y (n_1822));
AND2X1 g38943(.A (n_1227), .B (n_866), .Y (n_1519));
INVX1 g41951(.A (out_slt_127), .Y (n_217));
MX2X1 g29989(.A (n_322), .B (u0_slt9_r_170), .S0 (n_11319), .Y(n_11010));
MX2X1 g29988(.A (u1_sr_131), .B (in_slt_455), .S0 (out_le_184), .Y(n_11114));
MX2X1 g29987(.A (u1_sr_131), .B (in_slt_433), .S0 (out_le_183), .Y(n_11115));
MX2X1 g29986(.A (u1_sr_131), .B (in_slt_411), .S0 (out_le_182), .Y(n_11116));
MX2X1 g29985(.A (u1_sr_131), .B (in_slt_841), .S0 (out_le_181), .Y(n_11117));
MX2X1 g29984(.A (in_slt_742), .B (u1_sr_131), .S0 (out_le), .Y(n_11118));
INVX1 g42245(.A (out_slt_176), .Y (n_150));
INVX1 g41997(.A (out_slt_140), .Y (n_299));
INVX1 g41994(.A (crac_out_847), .Y (n_306));
INVX1 g41871(.A (out_slt_165), .Y (n_372));
INVX1 g43109(.A (out_slt_117), .Y (n_101));
MX2X1 g29796(.A (n_265), .B (u0_slt7_r_136), .S0 (n_11319), .Y(n_11249));
MX2X1 g29794(.A (n_375), .B (u0_slt7_r_137), .S0 (n_11389), .Y(n_11250));
MX2X1 g29792(.A (n_387), .B (u0_slt7_r_138), .S0 (n_11319), .Y(n_11251));
MX2X1 g29790(.A (n_229), .B (u0_slt7_r_139), .S0 (n_11389), .Y(n_11252));
MX2X1 g29798(.A (n_363), .B (u0_slt7_r_135), .S0 (n_11319), .Y(n_11248));
NOR3X1 g35841(.A (n_1213), .B (n_4076), .C (u2_cnt_b5_b ), .Y(n_4095));
INVX1 g42169(.A (out_slt_95), .Y (n_332));
INVX1 g42160(.A (out_slt_93), .Y (n_320));
INVX1 g42577(.A (crac_out), .Y (n_392));
INVX1 g42689(.A (out_slt_120), .Y (n_117));
NAND4X1 g37053(.A (n_3964), .B (n_701), .C (n_711), .D (n_2596), .Y(n_4000));
INVX1 g43049(.A (out_slt_76), .Y (n_157));
MX2X1 g30754(.A (u1_sr_127), .B (in_slt_753), .S0 (out_le_180), .Y(n_9764));
MX2X1 g30755(.A (u1_sr_127), .B (in_slt_837), .S0 (out_le_181), .Y(n_9763));
MX2X1 g30756(.A (u1_sr_127), .B (in_slt_407), .S0 (out_le_182), .Y(n_9762));
MX2X1 g30757(.A (u1_sr_127), .B (in_slt_429), .S0 (out_le_183), .Y(n_9761));
MX2X1 g30753(.A (in_slt_738), .B (u1_sr_127), .S0 (out_le), .Y(n_9765));
MX2X1 g30758(.A (u1_sr_127), .B (in_slt_451), .S0 (out_le_184), .Y(n_9760));
NOR2X1 g37052(.A (n_2602), .B (u2_cnt_b6_b ), .Y (n_2603));
INVX1 g42694(.A (out_slt_126), .Y (n_201));
MX2X1 g29854(.A (n_383), .B (u0_slt9_r_185), .S0 (n_11319), .Y(n_11217));
MX2X1 g29856(.A (n_19), .B (u0_slt9_r_184), .S0 (n_11319), .Y(n_11216));
MX2X1 g29850(.A (n_57), .B (u0_slt8_r), .S0 (n_11389), .Y (n_11219));
MX2X1 g29852(.A (n_273), .B (u0_slt9_r_186), .S0 (n_11389), .Y(n_11218));
MX2X1 g29858(.A (n_150), .B (u0_slt9_r_183), .S0 (n_7042), .Y(n_11215));
NAND2X1 g38953(.A (n_1253), .B (u2_cnt_b2_b ), .Y (n_1829));
INVX1 g42306(.A (out_slt_131), .Y (n_387));
MX2X1 g35367(.A (u1_sr), .B (in_slt3), .S0 (out_le_182), .Y (n_6731));
AND2X1 g29606(.A (u0_slt2_r_36), .B (n_11395), .Y (n_11368));
MX2X1 g29580(.A (n_338), .B (u0_slt2_r_49), .S0 (n_6710), .Y(n_11385));
INVX1 g42127(.A (out_slt_139), .Y (n_399));
MX2X1 g30134(.A (u1_sr_128), .B (in_slt_452), .S0 (out_le_184), .Y(n_9954));
MX2X1 g30136(.A (n_9952), .B (u0_slt9_r_169), .S0 (n_11319), .Y(n_9953));
MX2X1 g30131(.A (u1_sr_128), .B (in_slt_838), .S0 (out_le_181), .Y(n_9957));
MX2X1 g30132(.A (u1_sr_128), .B (in_slt_408), .S0 (out_le_182), .Y(n_9956));
MX2X1 g30133(.A (u1_sr_128), .B (in_slt_430), .S0 (out_le_183), .Y(n_9955));
AND2X1 g29698(.A (u0_slt5_r_107), .B (n_11395), .Y (n_11306));
MX2X1 g29878(.A (n_191), .B (u0_slt9_r_173), .S0 (n_6710), .Y(n_11204));
MX2X1 g29692(.A (n_397), .B (u0_slt5_r_110), .S0 (n_7042), .Y(n_11310));
MX2X1 g29690(.A (n_333), .B (u0_slt4_r), .S0 (n_7042), .Y (n_11311));
MX2X1 g29872(.A (n_308), .B (u0_slt9_r_176), .S0 (n_6710), .Y(n_11207));
MX2X1 g29870(.A (n_302), .B (u0_slt9_r_177), .S0 (n_6710), .Y(n_11209));
AND2X1 g41597(.A (n_1355), .B (n_1100), .Y (n_674));
NOR2X1 g36374(.A (n_1829), .B (n_698), .Y (n_2631));
XOR2X1 g36085(.A (u2_cnt_b3_b ), .B (n_1829), .Y (n_2629));
AND2X1 g29524(.A (u0_slt0_r_3), .B (n_7042), .Y (n_11423));
MX2X1 g29818(.A (n_240), .B (u0_slt8_r_164), .S0 (n_6710), .Y(n_11238));
MX2X1 g29810(.A (n_22), .B (u0_slt7_r), .S0 (n_11389), .Y (n_11242));
MX2X1 g29812(.A (n_184), .B (u0_slt8_r_167), .S0 (n_11319), .Y(n_11241));
MX2X1 g29814(.A (n_328), .B (u0_slt8_r_166), .S0 (n_11319), .Y(n_11240));
MX2X1 g29816(.A (n_86), .B (u0_slt8_r_165), .S0 (n_11395), .Y(n_11239));
INVX1 g42015(.A (crac_out_851), .Y (n_149));
AND2X1 g29718(.A (u0_slt5_r_97), .B (n_7042), .Y (n_11296));
AND2X1 g29716(.A (u0_slt5_r_98), .B (n_7042), .Y (n_11297));
AND2X1 g29714(.A (u0_slt5_r_99), .B (n_11395), .Y (n_11298));
AND2X1 g29712(.A (u0_slt5_r_100), .B (n_11395), .Y (n_11299));
AND2X1 g29710(.A (u0_slt5_r_101), .B (n_11395), .Y (n_11300));
INVX1 g43052(.A (out_slt_142), .Y (n_10983));
INVX1 g42693(.A (crac_out_854), .Y (n_112));
INVX1 g42470(.A (out_slt_135), .Y (n_186));
INVX1 g42476(.A (out_slt_151), .Y (n_181));
MX2X1 g35368(.A (u1_sr_118), .B (in_slt_398), .S0 (out_le_182), .Y(n_6730));
MX2X1 g35369(.A (u1_sr_119), .B (in_slt_399), .S0 (out_le_182), .Y(n_6729));
MX2X1 g35490(.A (u1_sr_120), .B (in_slt_830), .S0 (out_le_181), .Y(n_7144));
MX2X1 g35363(.A (u1_sr_121), .B (in_slt_423), .S0 (out_le_183), .Y(n_7362));
MX2X1 g35361(.A (u1_sr_120), .B (in_slt_400), .S0 (out_le_182), .Y(n_7156));
MX2X1 g35366(.A (u1_sr_121), .B (in_slt_747), .S0 (out_le_180), .Y(n_7359));
MX2X1 g35364(.A (u1_sr_121), .B (in_slt_445), .S0 (out_le_184), .Y(n_7361));
MX2X1 g35365(.A (u1_sr_121), .B (in_slt_831), .S0 (out_le_181), .Y(n_7360));
XOR2X1 g38469(.A (n_684), .B (n_1253), .Y (n_1552));
MX2X1 g29832(.A (n_167), .B (u0_slt8_r_157), .S0 (n_11389), .Y(n_11231));
MX2X1 g29830(.A (n_181), .B (u0_slt8_r_158), .S0 (n_11319), .Y(n_11232));
MX2X1 g29836(.A (n_376), .B (u0_slt8_r_155), .S0 (n_11389), .Y(n_11228));
MX2X1 g29834(.A (n_384), .B (u0_slt8_r_156), .S0 (n_11319), .Y(n_11230));
MX2X1 g29838(.A (n_362), .B (u0_slt8_r_154), .S0 (n_11319), .Y(n_11227));
AND2X1 g29526(.A (u0_slt0_r_2), .B (n_11395), .Y (n_11421));
NAND2X1 g29520(.A (u0_slt0_r_5), .B (n_7042), .Y (n_11425));
AND2X1 g29522(.A (u0_slt0_r_4), .B (n_11395), .Y (n_11424));
AND2X1 g29528(.A (u0_slt0_r_1), .B (n_7042), .Y (n_11420));
NAND2X1 g38946(.A (n_2377), .B (u2_cnt_b3_b ), .Y (n_3964));
INVX1 g38942(.A (n_1519), .Y (n_1520));
BUFX3 g35776(.A (n_6734), .Y (n_7042));
MX2X1 g35374(.A (u1_sr_119), .B (in_slt_421), .S0 (out_le_183), .Y(n_6725));
MX2X1 g35376(.A (u1_sr), .B (in_slt6), .S0 (out_le_184), .Y (n_6724));
MX2X1 g29738(.A (n_114), .B (u0_slt6_r_126), .S0 (n_11319), .Y(n_11286));
AND2X1 g29730(.A (u0_slt5_r), .B (n_11395), .Y (n_11290));
AND2X1 g29732(.A (u0_slt6_r_129), .B (n_11395), .Y (n_11289));
MX2X1 g29734(.A (n_102), .B (u0_slt6_r_128), .S0 (n_11319), .Y(n_11288));
NOR2X1 g41322(.A (n_688), .B (n_701), .Y (n_1138));
MX2X1 g31318(.A (u1_sr_126), .B (in_slt_450), .S0 (out_le_184), .Y(n_9618));
INVX1 g42670(.A (out_slt_137), .Y (n_254));
INVX1 g42412(.A (out_slt_132), .Y (n_229));
MX2X1 g29509(.A (out_slt_22), .B (u0_slt0_r_10), .S0 (n_11389), .Y(n_11433));
MX2X1 g29507(.A (out_slt_23), .B (u0_slt0_r_11), .S0 (n_11389), .Y(n_11434));
MX2X1 g29505(.A (out_slt_24), .B (u0_slt0_r_12), .S0 (n_11389), .Y(n_11435));
MX2X1 g29503(.A (out_slt_25), .B (u0_slt0_r_13), .S0 (n_11389), .Y(n_11436));
AOI21X1 g29501(.A0 (u0_slt0_r_14), .A1 (n_7042), .B0 (n_7013), .Y(n_11437));
NAND3X1 g29500(.A (n_11437), .B (n_7043), .C (n_11426), .Y (n_11438));
INVX1 g42086(.A (out_slt_125), .Y (n_335));
INVX1 g42332(.A (crac_out_852), .Y (n_357));
MX2X1 g29736(.A (n_117), .B (u0_slt6_r_127), .S0 (n_11389), .Y(n_11287));
MX2X1 g29756(.A (n_266), .B (u0_slt6_r_117), .S0 (n_11319), .Y(n_11273));
MX2X1 g29754(.A (n_264), .B (u0_slt6_r_118), .S0 (n_6710), .Y(n_11274));
MX2X1 g29758(.A (n_166), .B (u0_slt6_r_116), .S0 (n_6710), .Y(n_11272));
NAND3X1 g37196(.A (n_1782), .B (n_2571), .C (n_3995), .Y (n_3996));
AOI21X1 g37195(.A0 (n_2592), .A1 (n_2596), .B0 (n_702), .Y (n_2597));
INVX1 g42654(.A (out_slt_171), .Y (n_152));
INVX1 g42439(.A (out_slt_153), .Y (n_76));
NAND2X1 g29519(.A (n_11425), .B (n_11426), .Y (n_11427));
NOR2X1 g38990(.A (n_1773), .B (n_2377), .Y (n_2378));
AND2X1 g29568(.A (u0_slt1_r_16), .B (n_11395), .Y (n_11393));
AND2X1 g29560(.A (u0_slt1_r_20), .B (n_11395), .Y (n_11399));
AND2X1 g29562(.A (u0_slt1_r_19), .B (n_11395), .Y (n_11397));
AND2X1 g29564(.A (u0_slt1_r_18), .B (n_11395), .Y (n_11396));
AND2X1 g29566(.A (u0_slt1_r_17), .B (n_11395), .Y (n_11394));
MX2X1 g29958(.A (u1_sr_132), .B (in_slt_842), .S0 (out_le_181), .Y(n_11169));
MX2X1 g29959(.A (u1_sr_132), .B (in_slt_412), .S0 (out_le_182), .Y(n_11168));
MX2X1 g29776(.A (n_399), .B (u0_slt7_r_146), .S0 (n_11319), .Y(n_11260));
MX2X1 g29770(.A (n_21), .B (u0_slt6_r), .S0 (n_11319), .Y (n_11264));
MX2X1 g29772(.A (n_223), .B (u0_slt7_r_148), .S0 (n_11389), .Y(n_11263));
MX2X1 g34916(.A (n_120), .B (u0_slt9_r), .S0 (n_11319), .Y (n_8211));
XOR2X1 g36736(.A (u2_cnt_b5_b ), .B (n_1774), .Y (n_4826));
INVX1 g42184(.A (out_slt_144), .Y (n_182));
MX2X1 g35380(.A (u1_sr_120), .B (in_slt_444), .S0 (out_le_184), .Y(n_7154));
XOR2X1 g35381(.A (u2_cnt_b4_b ), .B (n_2632), .Y (n_5448));
MX2X1 g29897(.A (u1_sr_135), .B (in_slt_415), .S0 (out_le_182), .Y(n_11201));
MX2X1 g29896(.A (u1_sr_135), .B (in_slt_845), .S0 (out_le_181), .Y(n_11202));
MX2X1 g29899(.A (u1_sr_135), .B (in_slt_459), .S0 (out_le_184), .Y(n_11199));
INVX1 g42761(.A (n_866), .Y (n_687));
MX2X1 g29542(.A (crac_out_864), .B (u0_slt1_r_29), .S0 (n_7042), .Y(n_11411));
MX2X1 g29540(.A (crac_out_865), .B (u0_slt1_r_30), .S0 (n_7042), .Y(n_11413));
MX2X1 g29546(.A (crac_out_862), .B (u0_slt1_r_27), .S0 (n_11389), .Y(n_11409));
MX2X1 g29544(.A (crac_out_863), .B (u0_slt1_r_28), .S0 (n_7042), .Y(n_11410));
MX2X1 g29548(.A (crac_out_861), .B (u0_slt1_r_26), .S0 (n_11389), .Y(n_11408));
INVX1 g42444(.A (out_slt7), .Y (n_184));
INVX1 g41923(.A (out_slt_152), .Y (n_212));
INVX1 g42376(.A (out_slt_104), .Y (n_10785));
INVX1 g43021(.A (n_1773), .Y (n_688));
MX2X1 g29932(.A (u1_sr_133), .B (in_slt_843), .S0 (out_le_181), .Y(n_11187));
MX2X1 g29933(.A (u1_sr_133), .B (in_slt_413), .S0 (out_le_182), .Y(n_11186));
MX2X1 g29934(.A (u1_sr_133), .B (in_slt_435), .S0 (out_le_183), .Y(n_11185));
MX2X1 g29935(.A (u1_sr_133), .B (in_slt_457), .S0 (out_le_184), .Y(n_11184));
INVX1 g42619(.A (out_slt_91), .Y (n_391));
INVX1 g42968(.A (out_slt_82), .Y (n_16));
INVX1 g42617(.A (out_slt_130), .Y (n_375));
INVX1 g36752(.A (suspended_o), .Y (n_6057));
MX2X1 g34908(.A (u1_sr_122), .B (in_slt_424), .S0 (out_le_183), .Y(n_7511));
NOR2X1 g41402(.A (n_684), .B (n_698), .Y (n_1227));
MX2X1 g31824(.A (u1_sr_125), .B (in_slt_449), .S0 (out_le_184), .Y(n_9527));
NAND4X1 g37372(.A (n_2592), .B (n_1784), .C (n_701), .D (n_1773), .Y(n_2593));
INVX1 g41928(.A (out_slt_119), .Y (n_114));
INVX1 g42573(.A (out_slt_174), .Y (n_297));
INVX1 g42396(.A (out_slt_155), .Y (n_237));
INVX1 g42310(.A (out_slt_154), .Y (n_228));
MX2X1 g29914(.A (n_359), .B (u0_slt9_r_171), .S0 (n_11319), .Y(n_11188));
MX2X1 g29910(.A (u1_sr_134), .B (in_slt_844), .S0 (out_le_181), .Y(n_11198));
MX2X1 g29911(.A (u1_sr_134), .B (in_slt_414), .S0 (out_le_182), .Y(n_11197));
MX2X1 g29912(.A (u1_sr_134), .B (in_slt_436), .S0 (out_le_183), .Y(n_11196));
MX2X1 g29913(.A (u1_sr_134), .B (in_slt_458), .S0 (out_le_184), .Y(n_11195));
INVX1 g41849(.A (out_slt_147), .Y (n_362));
MX2X1 g29666(.A (n_330), .B (u0_slt4_r_84), .S0 (n_11319), .Y(n_11327));
MX2X1 g29664(.A (n_103), .B (u0_slt4_r_85), .S0 (n_6710), .Y(n_11328));
MX2X1 g29662(.A (n_243), .B (u0_slt4_r_86), .S0 (n_11319), .Y(n_11329));
MX2X1 g29660(.A (n_248), .B (u0_slt4_r_87), .S0 (n_11319), .Y(n_11330));
MX2X1 g29668(.A (n_332), .B (u0_slt4_r_83), .S0 (n_7042), .Y(n_11326));
INVX1 g42804(.A (out_slt_87), .Y (n_373));
INVX1 g42807(.A (crac_out_855), .Y (n_56));
INVX1 g42941(.A (out_slt_98), .Y (n_243));
INVX1 g42492(.A (out_slt_172), .Y (n_203));
INVX1 g41847(.A (out_slt_20), .Y (n_1372));
INVX1 g42569(.A (out_slt8), .Y (n_273));
NAND3X1 g37186(.A (n_1824), .B (n_684), .C (u2_cnt_b3_b ), .Y(n_4076));
MX2X1 g29586(.A (n_112), .B (u0_slt2_r_46), .S0 (n_11319), .Y(n_11381));
MX2X1 g29584(.A (n_56), .B (u0_slt2_r_47), .S0 (n_11319), .Y(n_11383));
MX2X1 g29582(.A (n_138), .B (u0_slt2_r_48), .S0 (n_11319), .Y(n_11384));
MX2X1 g29588(.A (n_231), .B (u0_slt2_r_45), .S0 (n_11319), .Y(n_11379));
NAND2X1 g41579(.A (n_687), .B (n_698), .Y (n_1114));
INVX1 g42005(.A (out_slt_133), .Y (n_401));
INVX1 g42004(.A (out_slt_19), .Y (n_1355));
INVX1 g43063(.A (out_slt_75), .Y (n_398));
MX2X1 g29640(.A (n_211), .B (u0_slt3_r_58), .S0 (n_11319), .Y(n_11346));
MX2X1 g29642(.A (n_200), .B (u0_slt3_r_57), .S0 (n_11319), .Y(n_11344));
MX2X1 g29644(.A (n_348), .B (u0_slt3_r_56), .S0 (n_11389), .Y(n_11342));
MX2X1 g29646(.A (n_10976), .B (u0_slt3_r_55), .S0 (n_11389), .Y(n_11341));
MX2X1 g29648(.A (n_10978), .B (u0_slt3_r_54), .S0 (n_11389), .Y(n_11339));
INVX1 g42829(.A (out_slt_92), .Y (n_394));
INVX1 g42927(.A (out_slt_114), .Y (n_84));
NOR2X1 g41356(.A (n_688), .B (n_687), .Y (n_1253));
INVX1 g42214(.A (out_slt_106), .Y (n_304));
MX2X1 g29840(.A (n_352), .B (u0_slt8_r_153), .S0 (n_11389), .Y(n_11225));
INVX1 g42026(.A (out_slt_124), .Y (n_10988));
MX2X1 g35362(.A (u1_sr_117), .B (in_slt_397), .S0 (out_le_182), .Y(n_6732));
INVX1 g42612(.A (out_slt_100), .Y (n_396));
INVX1 g41825(.A (out_slt_17), .Y (n_7017));
INVX1 g43085(.A (out_slt_160), .Y (n_120));
INVX1 g43082(.A (out_slt_85), .Y (n_10790));
AND2X1 g38822(.A (n_674), .B (n_1372), .Y (n_1087));
MX2X1 g29628(.A (n_157), .B (u0_slt3_r_64), .S0 (n_11319), .Y(n_11353));
MX2X1 g29622(.A (n_282), .B (u0_slt3_r_67), .S0 (n_11395), .Y(n_11356));
MX2X1 g29620(.A (n_281), .B (u0_slt3_r_68), .S0 (n_11395), .Y(n_11358));
MX2X1 g29626(.A (n_195), .B (u0_slt3_r_65), .S0 (n_7042), .Y(n_11354));
MX2X1 g29624(.A (n_267), .B (u0_slt3_r_66), .S0 (n_7042), .Y(n_11355));
INVX1 g42843(.A (out_slt_79), .Y (n_282));
NAND2X1 g36550(.A (n_1773), .B (n_6057), .Y (n_5822));
NAND2X1 g36551(.A (n_1928), .B (n_6057), .Y (n_5821));
NAND2X1 g36553(.A (n_1552), .B (n_6057), .Y (n_5820));
INVX1 g42443(.A (out_slt_116), .Y (n_261));
AOI21X1 g35675(.A0 (n_440), .A1 (n_679), .B0 (n_7042), .Y (n_7013));
INVX1 g41792(.A (out_slt_71), .Y (n_230));
INVX1 g42547(.A (out_slt_89), .Y (n_370));
INVX1 g42048(.A (out_slt_84), .Y (n_333));
INVX4 g35795(.A (n_7003), .Y (n_11319));
NAND3X1 g39825(.A (u2_cnt_b3_b ), .B (n_701), .C (n_456), .Y (n_1469));
MX2X1 g29604(.A (n_392), .B (u0_slt2_r_37), .S0 (n_11319), .Y(n_11370));
MX2X1 g29600(.A (n_306), .B (u0_slt2_r_39), .S0 (n_11319), .Y(n_11372));
MX2X1 g29602(.A (n_227), .B (u0_slt2_r_38), .S0 (n_11319), .Y(n_11371));
AND2X1 g29608(.A (u0_slt2_r_35), .B (n_7042), .Y (n_11366));
AND2X1 g39821(.A (u2_cnt_b4_b ), .B (n_3995), .Y (n_1784));
NAND2X1 g41258(.A (n_684), .B (n_687), .Y (n_2377));
NOR2X1 g41257(.A (out_slt_25), .B (out_slt_24), .Y (n_440));
INVX1 g41787(.A (out_slt_148), .Y (n_376));
MX2X1 g29752(.A (n_290), .B (u0_slt6_r_119), .S0 (n_11319), .Y(n_11276));
MX2X1 g29750(.A (n_287), .B (u0_slt6_r_120), .S0 (n_11389), .Y(n_11278));
NAND4X1 g35478(.A (n_2631), .B (u2_cnt_b5_b ), .C (u2_cnt_b6_b ), .D(u2_cnt_b4_b ), .Y (n_4103));
INVX1 g42527(.A (out_slt_70), .Y (n_211));
INVX1 g42524(.A (out_slt_22), .Y (n_1301));
INVX1 g42257(.A (out_slt_111), .Y (n_264));
INVX1 g42251(.A (out_slt_99), .Y (n_248));
INVX1 g42259(.A (out_slt_86), .Y (n_10788));
OR2X1 g35584(.A (n_7042), .B (n_7017), .Y (n_11426));
MX2X1 g33188(.A (u1_sr_124), .B (in_slt_426), .S0 (out_le_183), .Y(n_9354));
MX2X1 g33189(.A (u1_sr_124), .B (in_slt_448), .S0 (out_le_184), .Y(n_9353));
MX2X1 g33185(.A (u1_sr_124), .B (in_slt_750), .S0 (out_le_180), .Y(n_9357));
MX2X1 g33186(.A (u1_sr_124), .B (in_slt_834), .S0 (out_le_181), .Y(n_9356));
MX2X1 g33187(.A (u1_sr_124), .B (in_slt_404), .S0 (out_le_182), .Y(n_9355));
NAND2X1 g34715(.A (n_5448), .B (n_6057), .Y (n_6058));
NAND3X1 g36696(.A (n_1822), .B (n_1824), .C (u2_cnt_b2_b ), .Y(n_1823));
NOR2X1 g36695(.A (n_1785), .B (n_4076), .Y (n_4077));
INVX1 g42066(.A (out_slt_103), .Y (n_21));
AND2X1 g41660(.A (n_456), .B (n_711), .Y (n_3995));
INVX1 g42659(.A (out_slt_118), .Y (n_113));
NAND2X1 g33371(.A (n_5635), .B (n_6057), .Y (n_6066));
INVX1 g42656(.A (out_slt_107), .Y (n_262));
INVX1 g42500(.A (out_slt_150), .Y (n_167));
INVX1 g42504(.A (out_slt_97), .Y (n_103));
INVX1 g42506(.A (crac_out_853), .Y (n_231));
MX2X1 g30080(.A (u1_sr_129), .B (in_slt_431), .S0 (out_le_183), .Y(n_10802));
MX2X1 g30081(.A (u1_sr_129), .B (in_slt_453), .S0 (out_le_184), .Y(n_10800));
INVX1 g42212(.A (out_slt_112), .Y (n_290));
AND2X1 g41424(.A (n_1374), .B (n_1301), .Y (n_679));
INVX1 g42312(.A (out_slt_94), .Y (n_321));
MX2X1 g34080(.A (u1_sr_123), .B (in_slt_833), .S0 (out_le_181), .Y(n_8257));
MX2X1 g34081(.A (u1_sr_123), .B (in_slt_403), .S0 (out_le_182), .Y(n_8256));
MX2X1 g34082(.A (u1_sr_123), .B (in_slt_425), .S0 (out_le_183), .Y(n_8255));
MX2X1 g34083(.A (u1_sr_123), .B (in_slt_447), .S0 (out_le_184), .Y(n_8254));
INVX1 g42318(.A (out_slt_88), .Y (n_380));
OR2X1 g41218(.A (n_701), .B (n_711), .Y (n_702));
INVX1 g42777(.A (out_slt_69), .Y (n_200));
NOR2X1 g35633(.A (n_11395), .B (out_slt9), .Y (n_7231));
INVX1 g42299(.A (out_slt_177), .Y (n_19));
INVX1 g42295(.A (out_slt_134), .Y (n_259));
INVX1 g42236(.A (out_slt_141), .Y (n_57));
INVX1 g41985(.A (out_slt_163), .Y (n_322));
INVX1 g42237(.A (out_slt_90), .Y (n_351));
INVX1 g42179(.A (out_slt_149), .Y (n_384));
MX2X1 g29784(.A (n_186), .B (u0_slt7_r_142), .S0 (n_11319), .Y(n_11255));
MX2X1 g29786(.A (n_259), .B (u0_slt7_r_141), .S0 (n_11319), .Y(n_11254));
MX2X1 g29780(.A (n_254), .B (u0_slt7_r_144), .S0 (n_11389), .Y(n_11257));
MX2X1 g29782(.A (n_134), .B (u0_slt7_r_143), .S0 (n_11389), .Y(n_11256));
MX2X1 g29788(.A (n_401), .B (u0_slt7_r_140), .S0 (n_11389), .Y(n_11253));
INVX1 g42231(.A (out_slt_23), .Y (n_1374));
INVX1 g42177(.A (out_slt_68), .Y (n_348));
INVX1 g41980(.A (out_slt_109), .Y (n_166));
MX2X1 g29846(.A (n_10981), .B (u0_slt8_r_150), .S0 (n_11319), .Y(n_11221));
MX2X1 g29844(.A (n_182), .B (u0_slt8_r_151), .S0 (n_11389), .Y(n_11223));
MX2X1 g29842(.A (n_280), .B (u0_slt8_r_152), .S0 (n_11389), .Y(n_11224));
MX2X1 g29848(.A (n_10983), .B (u0_slt8_r_149), .S0 (n_11319), .Y(n_11220));
MX2X1 g29960(.A (u1_sr_132), .B (in_slt_434), .S0 (out_le_183), .Y(n_11167));
NAND4X1 g37007(.A (u2_cnt_b2_b ), .B (n_1138), .C (n_3995), .D(n_2596), .Y (n_2604));
NAND2X1 g35463(.A (n_2629), .B (n_6057), .Y (n_6052));
NAND3X1 g39719(.A (n_2596), .B (n_1212), .C (n_711), .Y (n_1213));

endmodule