
module buf1 (out, in);
    output out;
    input in;
    buf (out, in);
endmodule
    module clk_i_domain (scan_enable, scan_data_in, scan_data_out, clk_i, in_slt_434, in_slt_447, in_slt_450, in_slt_413, in_valid_8, wb_data_i_b6_b, n_290, n_287, n_84, in_slt_425, in_slt_426, wb_data_i_b21_b, in_slt_453, wb_data_i_b9_b, wb_data_i_b1_b, in_slt_742, wb_data_i_b13_b, in_slt_410, in_slt_411, in_slt_407, in_slt_431, in_slt_444, in_slt_456, n_7017, n_1100, in_slt_459, in_slt_457, in_slt_437, in_slt_435, dma_ack_i_b6_b, in_slt_458, in_slt_405, in_slt_399, in_slt_404, n_265, n_375, n_201, n_217, n_363, n_1557, wb_cyc_i, wb_stb_i, n_1559, wb_data_i_b30_b, n_82, n_19, n_383, wb_addr_i_b5_b, dma_ack_i_b8_b, in_slt_433, in_slt_443, wb_data_i_b22_b, in_slt_424, in_slt_420, in_slt_430, in_slt_406, n_182, n_228, n_237, n_86, n_240, n_328, in_slt_403, in_slt_739, in_slt_402, in_slt6, n_109, n_281, n_282, n_267, n_329, n_308, n_16, n_152, n_302, wb_data_i_b17_b, n_1355, n_793, n_1277, n_1553, wb_addr_i_b3_b, dma_ack_i_b3_b, dma_ack_i_b2_b, dma_ack_i_b1_b, dma_ack_i_b0_b, dma_ack_i_b5_b, dma_ack_i_b4_b, wb_data_i_b23_b, wb_data_i_b16_b, wb_addr_i_b6_b, wb_data_i_b3_b, in_slt_415, in_slt_397, in_slt_398, in_slt_446, wb_data_i_b15_b, wb_data_i_b24_b, in_slt_401, n_227, n_306, n_177, n_170, n_338, n_179, n_138, n_130, n_10790, n_10788, n_10785, n_10783, in_slt_409, n_9952, n_9602, n_10976, n_10978, n_10981, bit_clk_pad_i, in_slt_836, in_slt_455, wb_addr_i_b2_b, wb_data_i_b18_b, in_slt_412, in_slt_422, in_slt_408, in_slt_432, wb_addr_i_b31_b, wb_addr_i_b29_b, wb_data_i_b8_b, in_slt_436, in_slt_427, wb_data_i_b0_b, n_1374, n_370, n_380, n_391, n_351, n_361, n_373, n_394, in_slt_428, in_slt_449, in_slt_843, wb_data_i_b10_b, in_slt_830, in_slt_842, in_slt_840, n_6057, in_slt_423, in_slt_831, in_slt_429, wb_data_i_b31_b, in_slt_441, n_335, n_134, n_186, n_163, n_254, n_399, n_230, n_299, in_slt_445, in_slt_454, in_slt_448, n_1372, wb_data_i_b25_b, wb_data_i_b5_b, wb_addr_i_b4_b, n_113, n_101, n_261, n_300, n_102, n_117, n_114, n_304, in_slt_747, in_slt_414, in_slt_400, in_slt_442, in_slt_452, n_1301, wb_data_i_b28_b, in_slt_748, n_103, n_191, n_183, n_359, n_372, n_322, n_1233, n_212, n_181, n_167, n_243, n_332, n_76, wb_data_i_b27_b, dma_ack_i_b7_b, n_341, wb_data_i_b12_b, n_157, n_195, n_362, n_376, n_280, n_352, n_389, n_398, n_384, in_slt4, in_slt_738, wb_data_i_b2_b, in_slt_749, wb_data_i_b7_b, in_slt_451, n_348, n_297, n_200, n_208, n_203, n_263, n_150, n_211, in_slt3, wb_we_i, n_112, n_311, n_149, n_357, n_231, valid, in_slt_753, in_valid_9, in_slt_750, wb_data_i_b11_b, wb_data_i_b26_b, in_slt_421, n_392, n_10983, n_10988, wb_addr_i_b30_b, n_79, n_56, n_71, in_slt_844, in_slt_845, in_slt_838, in_valid, wb_data_i_b20_b, in_slt_752, wb_data_i_b29_b, wb_data_i_b14_b, in_slt_736, n_396, n_160, n_248, n_321, n_330, n_320, n_295, in_slt_833, wb_data_i_b4_b, wb_data_i_b19_b, in_slt_837, in_slt_841, in_slt_839, in_slt_832, in_slt_419, in_slt_834, n_10990, n_401, n_259, n_166, n_266, n_262, n_234, n_387, n_229, n_264, in_slt_835, wb_data_o_b27_b, wb_data_o_b20_b, wb_data_o_b28_b, out_slt_152, out_slt_161, out_slt_145, out_slt_164, out_slt_97, out_slt_85, out_slt_140, out_slt_116, wb_data_o_b16_b, out_slt_135, out_slt_121, out_slt_176, out_slt_173, out_slt_83, out_slt_115, out_slt_74, crac_out_860, out_slt_108, out_slt_124, out_slt_94, wb_data_o_b2_b, out_slt_91, out_slt_22, crac_out_847, out_slt_159, wb_data_o_b21_b, out_slt_151, wb_data_o_b29_b, out_slt_142, out_slt_132, out_slt_163, out_slt_119, out_slt_69, wb_data_o_b11_b, out_slt_66, out_slt_170, crac_out_850, out_slt_82, wb_data_o_b31_b, out_slt_105, crac_out_859, out_slt_102, out_slt_154, wb_data_o_b25_b, out_slt_123, out_slt_167, wb_data_o_b3_b, out_slt_99, out_slt_114, out_slt_133, wb_data_o_b14_b, out_slt_17, out_slt_178, out_slt_67, out_slt_77, wb_data_o_b30_b, crac_out_858, out_slt_106, out_slt_23, out_slt_126, out_slt_96, wb_data_o_b0_b, crac_out, out_slt_90, crac_out_854, wb_data_o_b9_b, out_slt_153, out_slt_144, out_slt_162, out_slt_138, out_slt_139, wb_data_o_b26_b, out_slt_117, out_slt_72, out_slt_71, wb_data_o_b17_b, out_slt_172, out_slt_175, out_slt_79, out_slt_76, out_slt_149, crac_out_857, wb_data_o_b6_b, out_slt_156, out_slt_19, wb_data_o_b23_b, out_slt_125, out_slt_93, out_slt_146, wb_data_o_b1_b, out_slt_92, out_slt_89, crac_out_846, out_slt_120, out_slt_112, out_slt_131, wb_data_o_b12_b, out_slt_68, out_slt_169, out_slt_78, crac_out_856, out_slt_129, out_slt_104, out_slt_128, out_slt_98, out_slt_88, crac_out_851, wb_data_o_b7_b, out_slt_155, out_slt_101, wb_data_o_b24_b, out_slt_168, out_slt_147, out_slt_136, out_slt_73, out_slt_70, wb_data_o_b15_b, out_slt_174, out_slt_177, out_slt_81, crac_out_848, out_slt_109, out_slt_110, crac_out_855, out_slt_158, out_slt_150, out_slt_127, out_slt_95, out_slt_143, out_slt_166, out_slt_148, out_slt_87, crac_out_853, crac_out_852, out_slt_118, wb_data_o_b19_b, out_slt_18, out_slt_137, wb_data_o_b10_b, out_slt_171, out_slt_80, int_o, out_slt_111, wb_data_o_b4_b, out_slt_100, out_slt_86, crac_out_849, wb_data_o_b5_b, out_slt_157, wb_data_o_b22_b, out_slt_134, out_slt_165, out_slt_20, wb_data_o_b8_b, out_slt_113, wb_data_o_b18_b, wb_data_o_b13_b, out_slt_75, out_slt_107);

input scan_enable, scan_data_in, clk_i, in_slt_434, in_slt_447, in_slt_450, in_slt_413, in_valid_8, wb_data_i_b6_b, n_290, n_287, n_84, in_slt_425, in_slt_426, wb_data_i_b21_b, in_slt_453, wb_data_i_b9_b, wb_data_i_b1_b, in_slt_742, wb_data_i_b13_b, in_slt_410, in_slt_411, in_slt_407, in_slt_431, in_slt_444, in_slt_456, n_7017, n_1100, in_slt_459, in_slt_457, in_slt_437, in_slt_435, dma_ack_i_b6_b, in_slt_458, in_slt_405, in_slt_399, in_slt_404, n_265, n_375, n_201, n_217, n_363, n_1557, wb_cyc_i, wb_stb_i, n_1559, wb_data_i_b30_b, n_82, n_19, n_383, wb_addr_i_b5_b, dma_ack_i_b8_b, in_slt_433, in_slt_443, wb_data_i_b22_b, in_slt_424, in_slt_420, in_slt_430, in_slt_406, n_182, n_228, n_237, n_86, n_240, n_328, in_slt_403, in_slt_739, in_slt_402, in_slt6, n_109, n_281, n_282, n_267, n_329, n_308, n_16, n_152, n_302, wb_data_i_b17_b, n_1355, n_793, n_1277, n_1553, wb_addr_i_b3_b, dma_ack_i_b3_b, dma_ack_i_b2_b, dma_ack_i_b1_b, dma_ack_i_b0_b, dma_ack_i_b5_b, dma_ack_i_b4_b, wb_data_i_b23_b, wb_data_i_b16_b, wb_addr_i_b6_b, wb_data_i_b3_b, in_slt_415, in_slt_397, in_slt_398, in_slt_446, wb_data_i_b15_b, wb_data_i_b24_b, in_slt_401, n_227, n_306, n_177, n_170, n_338, n_179, n_138, n_130, n_10790, n_10788, n_10785, n_10783, in_slt_409, n_9952, n_9602, n_10976, n_10978, n_10981, bit_clk_pad_i, in_slt_836, in_slt_455, wb_addr_i_b2_b, wb_data_i_b18_b, in_slt_412, in_slt_422, in_slt_408, in_slt_432, wb_addr_i_b31_b, wb_addr_i_b29_b, wb_data_i_b8_b, in_slt_436, in_slt_427, wb_data_i_b0_b, n_1374, n_370, n_380, n_391, n_351, n_361, n_373, n_394, in_slt_428, in_slt_449, in_slt_843, wb_data_i_b10_b, in_slt_830, in_slt_842, in_slt_840, n_6057, in_slt_423, in_slt_831, in_slt_429, wb_data_i_b31_b, in_slt_441, n_335, n_134, n_186, n_163, n_254, n_399, n_230, n_299, in_slt_445, in_slt_454, in_slt_448, n_1372, wb_data_i_b25_b, wb_data_i_b5_b, wb_addr_i_b4_b, n_113, n_101, n_261, n_300, n_102, n_117, n_114, n_304, in_slt_747, in_slt_414, in_slt_400, in_slt_442, in_slt_452, n_1301, wb_data_i_b28_b, in_slt_748, n_103, n_191, n_183, n_359, n_372, n_322, n_1233, n_212, n_181, n_167, n_243, n_332, n_76, wb_data_i_b27_b, dma_ack_i_b7_b, n_341, wb_data_i_b12_b, n_157, n_195, n_362, n_376, n_280, n_352, n_389, n_398, n_384, in_slt4, in_slt_738, wb_data_i_b2_b, in_slt_749, wb_data_i_b7_b, in_slt_451, n_348, n_297, n_200, n_208, n_203, n_263, n_150, n_211, in_slt3, wb_we_i, n_112, n_311, n_149, n_357, n_231, valid, in_slt_753, in_valid_9, in_slt_750, wb_data_i_b11_b, wb_data_i_b26_b, in_slt_421, n_392, n_10983, n_10988, wb_addr_i_b30_b, n_79, n_56, n_71, in_slt_844, in_slt_845, in_slt_838, in_valid, wb_data_i_b20_b, in_slt_752, wb_data_i_b29_b, wb_data_i_b14_b, in_slt_736, n_396, n_160, n_248, n_321, n_330, n_320, n_295, in_slt_833, wb_data_i_b4_b, wb_data_i_b19_b, in_slt_837, in_slt_841, in_slt_839, in_slt_832, in_slt_419, in_slt_834, n_10990, n_401, n_259, n_166, n_266, n_262, n_234, n_387, n_229, n_264, in_slt_835;
output scan_data_out, wb_data_o_b27_b, wb_data_o_b20_b, wb_data_o_b28_b, out_slt_152, out_slt_161, out_slt_145, out_slt_164, out_slt_97, out_slt_85, out_slt_140, out_slt_116, wb_data_o_b16_b, out_slt_135, out_slt_121, out_slt_176, out_slt_173, out_slt_83, out_slt_115, out_slt_74, crac_out_860, out_slt_108, out_slt_124, out_slt_94, wb_data_o_b2_b, out_slt_91, out_slt_22, crac_out_847, out_slt_159, wb_data_o_b21_b, out_slt_151, wb_data_o_b29_b, out_slt_142, out_slt_132, out_slt_163, out_slt_119, out_slt_69, wb_data_o_b11_b, out_slt_66, out_slt_170, crac_out_850, out_slt_82, wb_data_o_b31_b, out_slt_105, crac_out_859, out_slt_102, out_slt_154, wb_data_o_b25_b, out_slt_123, out_slt_167, wb_data_o_b3_b, out_slt_99, out_slt_114, out_slt_133, wb_data_o_b14_b, out_slt_17, out_slt_178, out_slt_67, out_slt_77, wb_data_o_b30_b, crac_out_858, out_slt_106, out_slt_23, out_slt_126, out_slt_96, wb_data_o_b0_b, crac_out, out_slt_90, crac_out_854, wb_data_o_b9_b, out_slt_153, out_slt_144, out_slt_162, out_slt_138, out_slt_139, wb_data_o_b26_b, out_slt_117, out_slt_72, out_slt_71, wb_data_o_b17_b, out_slt_172, out_slt_175, out_slt_79, out_slt_76, out_slt_149, crac_out_857, wb_data_o_b6_b, out_slt_156, out_slt_19, wb_data_o_b23_b, out_slt_125, out_slt_93, out_slt_146, wb_data_o_b1_b, out_slt_92, out_slt_89, crac_out_846, out_slt_120, out_slt_112, out_slt_131, wb_data_o_b12_b, out_slt_68, out_slt_169, out_slt_78, crac_out_856, out_slt_129, out_slt_104, out_slt_128, out_slt_98, out_slt_88, crac_out_851, wb_data_o_b7_b, out_slt_155, out_slt_101, wb_data_o_b24_b, out_slt_168, out_slt_147, out_slt_136, out_slt_73, out_slt_70, wb_data_o_b15_b, out_slt_174, out_slt_177, out_slt_81, crac_out_848, out_slt_109, out_slt_110, crac_out_855, out_slt_158, out_slt_150, out_slt_127, out_slt_95, out_slt_143, out_slt_166, out_slt_148, out_slt_87, crac_out_853, crac_out_852, out_slt_118, wb_data_o_b19_b, out_slt_18, out_slt_137, wb_data_o_b10_b, out_slt_171, out_slt_80, int_o, out_slt_111, wb_data_o_b4_b, out_slt_100, out_slt_86, crac_out_849, wb_data_o_b5_b, out_slt_157, wb_data_o_b22_b, out_slt_134, out_slt_165, out_slt_20, wb_data_o_b8_b, out_slt_113, wb_data_o_b18_b, wb_data_o_b13_b, out_slt_75, out_slt_107;
wire n_8047;
wire u8_mem_b3_b_122;
wire n_7976;
wire n_716;
wire n_715;
wire u15_rdd3;
wire n_10349;
wire n_5502;
wire n_10376;
wire n_8046;
wire u4_mem_b1_b_75;
wire n_7984;
wire n_2864;
wire wb_din_690;
wire n_4599;
wire n_3264;
wire n_2889;
wire n_1675;
wire n_379;
wire n_2544;
wire n_5359;
wire n_1316;
wire n_3917;
wire n_2404;
wire n_2250;
wire n_1678;
wire n_2558;
wire n_1677;
wire n_1676;
wire n_1839;
wire n_1681;
wire n_2502;
wire n_1680;
wire n_1679;
wire n_1859;
wire n_2548;
wire n_147;
wire n_940;
wire n_5512;
wire n_2551;
wire n_2550;
wire n_2549;
wire n_2534;
wire n_5215;
wire n_1523;
wire n_4234;
wire n_3916;
wire n_2444;
wire n_2320;
wire n_2628;
wire n_143;
wire n_2530;
wire n_2627;
wire n_11974;
wire n_7251;
wire n_7188;
wire n_10518;
wire n_11990;
wire n_7314;
wire n_7094;
wire n_11954;
wire n_7253;
wire n_7016;
wire n_11978;
wire n_7315;
wire n_7189;
wire n_11952;
wire n_7316;
wire n_6918;
wire n_11968;
wire n_7254;
wire n_7190;
wire n_11970;
wire n_7255;
wire n_7192;
wire n_11964;
wire n_7257;
wire n_7193;
wire n_4788;
wire u9_mem_b1_b_143;
wire n_4755;
wire n_4783;
wire n_4789;
wire u9_mem_b1_b_141;
wire n_4757;
wire n_4785;
wire u9_mem_b1_b_146;
wire n_4772;
wire u7_mem_b2_b_55;
wire n_8998;
wire n_4782;
wire u9_mem_b1_b_148;
wire n_4764;
wire n_4784;
wire u9_mem_b1_b_147;
wire n_4769;
wire n_11972;
wire n_7249;
wire n_7186;
wire n_10523;
wire n_7250;
wire n_7093;
wire u3_mem_b2_b_53;
wire n_9071;
wire n_742;
wire n_1819;
wire u5_mem_b0_b_93;
wire n_8786;
wire ic0_int_set_719;
wire n_7364;
wire u4_mem_b2_b_36;
wire n_8267;
wire n_8568;
wire wb_din_672;
wire n_8567;
wire n_8538;
wire n_8051;
wire u4_mem_b1_b_72;
wire u5_mem_b1_b_62;
wire n_9282;
wire u10_mem_b1_b_125;
wire n_10180;
wire n_8560;
wire wb_din_677;
wire oc2_cfg_984;
wire n_1441;
wire u26_ps_cnt_b1_b;
wire n_529;
wire n_819;
wire n_858;
wire n_627;
wire n_626;
wire n_1929;
wire u8_wp_b1_b;
wire n_12280;
wire n_6350;
wire n_6349;
wire n_6486;
wire n_6359;
wire n_6348;
wire n_6347;
wire n_6547;
wire n_6354;
wire n_6353;
wire n_6442;
wire n_6352;
wire n_6351;
wire n_6544;
wire n_6358;
wire n_6357;
wire n_6497;
wire n_6356;
wire n_6355;
wire n_6444;
wire u11_mem_b0_b_162;
wire n_10817;
wire n_5950;
wire n_5949;
wire n_6008;
wire n_6341;
wire n_1333;
wire u5_mem_b3_b_136;
wire n_1543;
wire u12_we2;
wire n_870;
wire n_6345;
wire n_6344;
wire n_6483;
wire n_5948;
wire n_5947;
wire n_5983;
wire n_39;
wire u10_mem_b2_b_108;
wire n_3502;
wire n_12826;
wire u3_mem_b0_b_108;
wire n_6942;
wire u9_mem_b1_b_124;
wire n_11043;
wire n_862;
wire n_1447;
wire n_494;
wire n_1446;
wire u8_rp_b3_b;
wire u8_wp_b2_b;
wire n_7328;
wire n_6818;
wire n_6135;
wire n_12145;
wire n_7278;
wire n_6313;
wire n_6133;
wire n_7324;
wire n_9605;
wire n_9604;
wire n_9554;
wire n_1208;
wire n_7160;
wire n_9503;
wire n_9553;
wire n_9552;
wire n_1071;
wire n_7036;
wire n_9560;
wire n_9551;
wire n_9550;
wire n_1130;
wire n_7035;
wire n_9501;
wire n_8848;
wire n_8847;
wire n_7532;
wire n_7527;
wire n_1116;
wire n_7034;
wire n_9499;
wire n_9445;
wire n_9444;
wire n_8208;
wire n_8206;
wire n_8844;
wire n_8843;
wire n_7529;
wire n_7525;
wire n_11934;
wire n_12357;
wire n_3509;
wire u6_mem_b2_b_45;
wire n_3474;
wire n_7108;
wire n_2583;
wire n_4716;
wire n_7353;
wire n_7107;
wire n_4665;
wire n_7151;
wire n_4662;
wire n_4105;
wire n_1292;
wire n_4104;
wire n_6708;
wire n_877;
wire n_1221;
wire i3_re;
wire n_6707;
wire n_1232;
wire n_2364;
wire i4_re;
wire n_11095;
wire n_11965;
wire n_11086;
wire n_11094;
wire n_11971;
wire n_5827;
wire n_10909;
wire n_9915;
wire n_9798;
wire n_10916;
wire n_10908;
wire n_9914;
wire n_9797;
wire n_2485;
wire n_10911;
wire n_12813;
wire n_12814;
wire n_10910;
wire n_12815;
wire n_12816;
wire n_10913;
wire n_12610;
wire n_11999;
wire n_10921;
wire n_10912;
wire n_12811;
wire n_12812;
wire n_10996;
wire n_10786;
wire n_10994;
wire n_10995;
wire n_10784;
wire n_12385;
wire n_12384;
wire n_2513;
wire n_1040;
wire n_12389;
wire n_4080;
wire n_1068;
wire u7_rp_b3_b;
wire n_5702;
wire n_6226;
wire i3_dout_587;
wire n_4051;
wire n_3575;
wire u3_mem_b0_b_94;
wire wb_din_664;
wire n_3807;
wire n_11712;
wire u6_mem_b1_b_64;
wire n_4253;
wire n_3572;
wire u3_mem_b0_b_98;
wire wb_din_668;
wire n_6715;
wire n_1080;
wire i6_re;
wire n_11461;
wire n_11798;
wire u8_mem_b0_b_105;
wire n_3573;
wire u6_mem_b0_b_109;
wire wb_din_679;
wire n_3632;
wire n_7140;
wire n_5592;
wire n_4731;
wire n_4192;
wire u4_mem_b1_b_61;
wire n_12259;
wire n_11714;
wire u6_mem_b1_b_65;
wire n_12169;
wire n_3571;
wire u7_mem_b0_b_115;
wire wb_din_685;
wire n_3622;
wire n_4128;
wire u7_mem_b2_b_52;
wire n_12650;
wire n_2964;
wire n_3332;
wire n_2801;
wire u10_mem_b3_b_58;
wire n_10567;
wire i4_dout_599;
wire n_4022;
wire n_2969;
wire u7_mem_b2_b_35;
wire n_12654;
wire n_4751;
wire n_2302;
wire n_3569;
wire u7_mem_b0_b_113;
wire wb_din_683;
wire n_2249;
wire n_2325;
wire n_4129;
wire u7_mem_b2_b_51;
wire n_12645;
wire n_2965;
wire n_4996;
wire n_2720;
wire n_2966;
wire u7_mem_b2_b_37;
wire n_3567;
wire u6_mem_b0_b_104;
wire wb_din_674;
wire i6_dout_654;
wire n_4010;
wire n_3188;
wire u7_mem_b2_b_38;
wire n_12641;
wire n_4560;
wire n_1360;
wire n_10542;
wire n_6481;
wire n_419;
wire n_10513;
wire n_10543;
wire n_5985;
wire n_5984;
wire n_10215;
wire n_6477;
wire n_6476;
wire n_10315;
wire n_10540;
wire n_6480;
wire n_6479;
wire n_10537;
wire n_10546;
wire n_6549;
wire n_6548;
wire n_10547;
wire n_6488;
wire n_6487;
wire n_10544;
wire n_5982;
wire n_5981;
wire n_10565;
wire n_10545;
wire n_6485;
wire n_6484;
wire n_10214;
wire n_6469;
wire n_6468;
wire n_10539;
wire n_6474;
wire n_433;
wire n_2440;
wire u6_mem_b3_b_147;
wire n_2465;
wire u11_mem_b3_b_72;
wire n_10836;
wire n_5751;
wire n_5190;
wire n_5189;
wire n_634;
wire n_8730;
wire u7_mem_b0_b_93;
wire n_3616;
wire n_7493;
wire n_9393;
wire u7_mem_b0_b_121;
wire n_3635;
wire n_8733;
wire u7_mem_b0_b_119;
wire n_3610;
wire n_8735;
wire u7_mem_b0_b_118;
wire n_3636;
wire n_8731;
wire u7_mem_b0_b_120;
wire n_3613;
wire n_8732;
wire u7_mem_b0_b_92;
wire n_3612;
wire n_8738;
wire n_9394;
wire u7_mem_b0_b_114;
wire n_3639;
wire n_8736;
wire u7_mem_b0_b_117;
wire n_3607;
wire n_8737;
wire u7_mem_b0_b_116;
wire n_3638;
wire u9_mem_b2_b_100;
wire n_10284;
wire n_7136;
wire n_5589;
wire n_4724;
wire n_5315;
wire n_5920;
wire n_6821;
wire n_5844;
wire n_3460;
wire n_11804;
wire u8_mem_b0_b_113;
wire n_12806;
wire u5_mem_b2_b_42;
wire n_12823;
wire n_1501;
wire n_2691;
wire n_1488;
wire n_3463;
wire n_3089;
wire n_3008;
wire n_3465;
wire n_5138;
wire n_2702;
wire n_3466;
wire n_3415;
wire n_2618;
wire n_2617;
wire n_3944;
wire u13_ints_r_b22_b;
wire n_6749;
wire n_11451;
wire u8_mem_b0_b_100;
wire n_9325;
wire n_5072;
wire n_9349;
wire n_7955;
wire n_9327;
wire n_5074;
wire n_9326;
wire n_7956;
wire n_9328;
wire n_5075;
wire n_7958;
wire n_9329;
wire n_5077;
wire n_9336;
wire n_7959;
wire u11_din_tmp_51;
wire n_10114;
wire n_9331;
wire n_5080;
wire n_9333;
wire n_7961;
wire n_9332;
wire n_5081;
wire n_7962;
wire n_9334;
wire n_5082;
wire n_7963;
wire n_2695;
wire n_2780;
wire n_2729;
wire n_5922;
wire n_5851;
wire n_9322;
wire n_5068;
wire n_7953;
wire n_9324;
wire n_5071;
wire n_7954;
wire n_9009;
wire n_4466;
wire n_9055;
wire n_7675;
wire n_9011;
wire n_4314;
wire n_9010;
wire n_7676;
wire n_5923;
wire n_5853;
wire n_9019;
wire n_4406;
wire n_9043;
wire n_7683;
wire n_9020;
wire n_4404;
wire n_9034;
wire n_7684;
wire n_9016;
wire n_4424;
wire n_7681;
wire n_9018;
wire n_4318;
wire n_7682;
wire n_9014;
wire n_4316;
wire n_7679;
wire n_9015;
wire n_4317;
wire n_7680;
wire n_9012;
wire n_4452;
wire n_7677;
wire n_9013;
wire n_4315;
wire n_9038;
wire n_7678;
wire n_4777;
wire u9_mem_b2_b_109;
wire n_4776;
wire n_5732;
wire n_9161;
wire n_7428;
wire n_4779;
wire u9_mem_b2_b_107;
wire n_4778;
wire n_6898;
wire in_valid_s_1;
wire u3_mem_b0_b_97;
wire n_8249;
wire n_1480;
wire n_2712;
wire u5_mem_b0_b_100;
wire n_8808;
wire u13_intm_r_b21_b;
wire n_8507;
wire n_1660;
wire n_1756;
wire n_6360;
wire n_6503;
wire n_1643;
wire wb_din_666;
wire n_2412;
wire n_393;
wire ic0_cfg_1029;
wire n_8579;
wire n_8341;
wire n_2410;
wire u8_mem_b3_b_149;
wire n_2468;
wire n_4786;
wire u9_mem_b1_b_145;
wire n_4743;
wire u3_mem_b1_b_67;
wire n_8441;
wire n_2408;
wire u5_mem_b3_b_122;
wire n_3543;
wire n_2409;
wire u3_mem_b3_b_141;
wire n_2463;
wire n_4780;
wire u10_mem_b1_b_145;
wire n_4759;
wire n_5407;
wire n_11076;
wire n_7454;
wire n_4781;
wire u9_mem_b1_b_149;
wire n_4767;
wire n_5730;
wire u5_mem_b3_b_143;
wire n_9219;
wire i4_dout_618;
wire n_4037;
wire n_9750;
wire u11_wp_b0_b;
wire n_9631;
wire n_10949;
wire n_9931;
wire n_9833;
wire n_9933;
wire n_9751;
wire u10_wp_b3_b;
wire n_9564;
wire n_11823;
wire n_11827;
wire n_12638;
wire n_12636;
wire n_12634;
wire n_5818;
wire n_10103;
wire n_9932;
wire n_9930;
wire n_12659;
wire n_5442;
wire u11_rp_b0_b;
wire u11_wp_b1_b;
wire n_916;
wire n_5622;
wire n_1198;
wire u8_wp_b0_b;
wire n_1206;
wire n_5420;
wire n_1207;
wire n_6049;
wire n_1419;
wire n_1923;
wire n_1290;
wire u10_rp_b2_b;
wire n_514;
wire n_5616;
wire n_1421;
wire n_1921;
wire n_822;
wire u3_rp_b3_b;
wire u3_wp_b2_b;
wire n_477;
wire n_1926;
wire n_6841;
wire n_907;
wire u11_rp_b2_b;
wire u11_wp_b3_b;
wire n_522;
wire n_3577;
wire u3_mem_b0_b_121;
wire wb_din_691;
wire n_3576;
wire u6_mem_b0_b_107;
wire n_1025;
wire n_695;
wire n_5143;
wire u3_mem_b1_b_72;
wire n_5148;
wire n_2677;
wire n_6211;
wire n_4127;
wire n_2294;
wire n_3120;
wire n_1530;
wire n_5690;
wire n_6233;
wire n_4173;
wire n_2959;
wire n_3093;
wire n_1537;
wire n_6186;
wire n_3489;
wire n_2898;
wire n_2405;
wire n_5545;
wire n_5544;
wire n_3886;
wire u8_mem_b3_b;
wire n_3879;
wire n_1503;
wire n_3105;
wire n_2493;
wire n_1526;
wire n_5691;
wire u13_intm_r_b26_b;
wire n_8500;
wire n_6335;
wire u10_mem_b0_b_154;
wire n_6138;
wire n_4576;
wire n_5203;
wire n_784;
wire n_5795;
wire n_5252;
wire n_3980;
wire n_6823;
wire n_6779;
wire n_5924;
wire n_5855;
wire n_5925;
wire n_5833;
wire n_5926;
wire n_5835;
wire n_6825;
wire n_12746;
wire n_6824;
wire n_6309;
wire n_6237;
wire n_5248;
wire n_1284;
wire u12_we1;
wire n_6312;
wire n_6252;
wire n_5796;
wire n_5185;
wire n_5184;
wire u3_mem_b1_b_84;
wire n_8857;
wire n_12405;
wire n_1546;
wire u7_mem_b3_b_140;
wire n_12244;
wire n_12400;
wire u5_rp_b1_b;
wire n_12399;
wire n_12581;
wire n_12401;
wire n_12404;
wire n_2491;
wire u7_mem_b0_b_109;
wire n_12403;
wire n_4225;
wire u7_mem_b1_b_78;
wire n_12411;
wire n_12410;
wire n_1033;
wire u3_mem_b1_b_60;
wire n_8356;
wire n_3058;
wire n_3117;
wire n_2686;
wire out_slt7;
wire n_11111;
wire n_7485;
wire wb_din_689;
wire u5_mem_b2_b_39;
wire n_9272;
wire n_1516;
wire u7_mem_b3_b_141;
wire u4_mem_b3_b_151;
wire u6_mem_b2_b_55;
wire n_9127;
wire n_1694;
wire n_6900;
wire n_1835;
wire n_1693;
wire n_6849;
wire n_6886;
wire n_1760;
wire n_4607;
wire n_3531;
wire n_3367;
wire n_5219;
wire n_4140;
wire n_3366;
wire n_1692;
wire n_6033;
wire n_6013;
wire u8_mem_b1_b_83;
wire n_8920;
wire n_5218;
wire n_4219;
wire n_3362;
wire n_4078;
wire n_6030;
wire n_2553;
wire n_2365;
wire n_1249;
wire n_5955;
wire n_6010;
wire n_12252;
wire n_12258;
wire n_7453;
wire u6_mem_b1_b_89;
wire n_9160;
wire n_11073;
wire n_686;
wire n_685;
wire n_708;
wire n_9611;
wire n_8550;
wire oc2_cfg_987;
wire u3_mem_b0_b_113;
wire n_8701;
wire n_1064;
wire u10_wp_b1_b;
wire u10_wp_b2_b;
wire n_513;
wire u13_ints_r_b27_b;
wire ic2_int_set_723;
wire u7_rp_b0_b;
wire n_9871;
wire u10_din_tmp_44;
wire n_9860;
wire n_9869;
wire u10_din_tmp_45;
wire n_10364;
wire n_298;
wire n_10363;
wire n_236;
wire n_1968;
wire n_2144;
wire n_2755;
wire n_10369;
wire n_279;
wire n_9989;
wire n_11890;
wire n_1184;
wire n_10371;
wire n_81;
wire n_10385;
wire n_10370;
wire n_1627;
wire n_10365;
wire n_270;
wire n_10118;
wire n_5963;
wire n_5962;
wire n_10137;
wire n_10810;
wire n_9901;
wire n_10366;
wire n_275;
wire n_5175;
wire n_2867;
wire n_2876;
wire n_5174;
wire n_1812;
wire n_3442;
wire n_3892;
wire n_6457;
wire n_6591;
wire n_5178;
wire n_3419;
wire n_5180;
wire n_3003;
wire n_3429;
wire n_5179;
wire n_2396;
wire n_2844;
wire n_5176;
wire n_2852;
wire n_3160;
wire n_4552;
wire n_2383;
wire n_2301;
wire n_5177;
wire n_2375;
wire n_2891;
wire n_2503;
wire n_6394;
wire n_6537;
wire n_9795;
wire u15_rdd1;
wire n_9688;
wire n_9794;
wire crac_wr;
wire n_9689;
wire u7_wp_b1_b;
wire n_9455;
wire n_9571;
wire n_8210;
wire u14_u8_en_out_l2;
wire u5_mem_b1_b_81;
wire n_3239;
wire u11_mem_b3_b_65;
wire n_10654;
wire u10_mem_b2_b_97;
wire n_10325;
wire n_9712;
wire n_9711;
wire n_294;
wire n_8179;
wire n_991;
wire n_614;
wire n_7522;
wire n_7521;
wire wb_din_661;
wire n_6431;
wire u11_mem_b2_b_95;
wire n_1272;
wire n_12637;
wire n_12635;
wire n_11130;
wire n_6005;
wire u10_mem_b3_b;
wire u11_mem_b0_b_153;
wire n_10424;
wire n_6854;
wire u9_mem_b0_b_153;
wire u7_mem_b1_b_60;
wire n_9049;
wire wb_din_681;
wire n_11698;
wire u6_mem_b2_b_40;
wire n_11061;
wire n_6651;
wire n_6650;
wire n_6649;
wire n_6653;
wire n_6652;
wire n_6579;
wire n_5341;
wire n_6943;
wire n_6899;
wire n_6946;
wire n_6945;
wire n_6913;
wire n_6938;
wire n_6937;
wire n_6906;
wire n_6941;
wire n_6940;
wire n_6927;
wire n_6645;
wire n_6644;
wire n_6618;
wire u11_mem_b3_b_75;
wire n_10857;
wire n_6639;
wire n_6638;
wire n_6637;
wire n_6642;
wire n_6641;
wire n_6533;
wire n_1051;
wire n_704;
wire u2_to_cnt_b1_b;
wire n_11742;
wire u8_mem_b0_b_91;
wire n_3890;
wire u8_mem_b0_b_108;
wire n_2227;
wire n_2851;
wire n_2741;
wire n_2850;
wire u8_mem_b1_b_77;
wire n_12291;
wire n_12087;
wire n_12076;
wire i4_dout_619;
wire n_4818;
wire ic2_cfg_1045;
wire n_8604;
wire n_12079;
wire u8_mem_b2_b_29;
wire n_8871;
wire n_8930;
wire n_7396;
wire n_8433;
wire n_8449;
wire n_8453;
wire n_8457;
wire n_8464;
wire n_8438;
wire n_7612;
wire u8_mem_b1_b_73;
wire n_7611;
wire u8_mem_b1_b_74;
wire n_7614;
wire u8_mem_b1_b_70;
wire n_7613;
wire u8_mem_b1_b_72;
wire n_7608;
wire n_7607;
wire u3_mem_b1_b_90;
wire n_8101;
wire n_7610;
wire u8_mem_b1_b_76;
wire n_7609;
wire u8_mem_b3_b_133;
wire n_7606;
wire u8_mem_b1_b_78;
wire n_7605;
wire u8_mem_b1_b_79;
wire n_12631;
wire n_11855;
wire n_11020;
wire n_11142;
wire n_6839;
wire n_11136;
wire n_10960;
wire n_11526;
wire n_6836;
wire n_12589;
wire n_10963;
wire n_9753;
wire n_9581;
wire n_9650;
wire n_599;
wire n_9754;
wire n_9582;
wire n_9653;
wire n_690;
wire n_11505;
wire n_6059;
wire n_10959;
wire n_7455;
wire n_7301;
wire n_6696;
wire n_11522;
wire n_6842;
wire n_11126;
wire n_11005;
wire n_11520;
wire n_7049;
wire n_11131;
wire n_11007;
wire n_3256;
wire n_3255;
wire u5_mem_b0_b_97;
wire n_2321;
wire n_2330;
wire u7_mem_b0_b_91;
wire n_10970;
wire n_6756;
wire n_10328;
wire n_10985;
wire n_10971;
wire n_7010;
wire n_10330;
wire n_10992;
wire n_7475;
wire i4_dout;
wire n_7468;
wire n_7352;
wire n_6054;
wire n_5445;
wire u2_bit_clk_e;
wire u11_mem_b3_b_57;
wire n_10455;
wire u7_mem_b2_b_50;
wire n_9003;
wire n_6147;
wire n_3161;
wire n_2247;
wire n_3514;
wire n_1521;
wire n_10942;
wire u5_mem_b2_b_37;
wire n_9238;
wire n_4004;
wire n_1574;
wire n_1573;
wire n_5553;
wire n_11717;
wire n_11718;
wire n_2286;
wire n_2428;
wire n_6076;
wire n_12171;
wire n_4005;
wire n_1577;
wire n_1576;
wire n_5554;
wire u10_mem_b0_b_180;
wire n_10126;
wire n_11528;
wire n_9476;
wire u8_mem_b2_b_41;
wire n_8882;
wire u13_intm_r_b0_b;
wire n_8521;
wire u3_mem_b2_b_59;
wire n_8398;
wire n_10081;
wire n_9724;
wire n_9676;
wire n_9632;
wire n_9829;
wire wb_din_669;
wire n_4200;
wire u4_mem_b1_b_82;
wire n_12267;
wire u13_intm_r_b14_b;
wire n_8515;
wire n_2170;
wire n_2169;
wire n_2681;
wire u8_mem_b0_b_93;
wire n_8691;
wire n_8526;
wire n_8527;
wire n_2168;
wire n_2038;
wire n_2786;
wire u5_mem_b3_b_138;
wire n_9227;
wire u11_mem_b2_b_92;
wire n_10494;
wire n_8085;
wire u3_mem_b3_b_147;
wire n_8141;
wire n_8386;
wire n_4871;
wire n_9022;
wire n_8100;
wire n_8385;
wire n_4889;
wire n_8383;
wire n_8099;
wire n_8384;
wire n_5139;
wire n_8098;
wire u7_mem_b2_b_45;
wire n_8244;
wire n_6675;
wire n_7459;
wire n_8379;
wire n_5136;
wire n_8380;
wire n_8094;
wire n_8378;
wire n_5135;
wire n_8093;
wire n_8377;
wire n_4910;
wire n_8375;
wire n_8092;
wire ic1_cfg_1036;
wire n_8620;
wire n_10999;
wire u5_mem_b2_b_53;
wire n_9254;
wire n_5534;
wire n_5898;
wire n_7777;
wire u6_mem_b2_b_51;
wire n_7758;
wire n_8855;
wire n_4434;
wire n_7977;
wire n_7779;
wire u6_mem_b2_b_49;
wire n_7778;
wire u6_mem_b2_b_50;
wire u8_mem_b3_b_126;
wire n_8420;
wire n_3268;
wire u5_mem_b0_b_96;
wire n_7780;
wire u6_mem_b2_b_48;
wire n_11082;
wire u11_mem_b2_b_117;
wire n_10860;
wire n_8862;
wire n_4304;
wire n_8891;
wire n_7662;
wire n_8866;
wire n_4860;
wire n_8856;
wire n_7570;
wire n_8865;
wire n_4298;
wire n_8868;
wire n_7700;
wire n_5055;
wire u6_mem_b3_b_145;
wire n_5059;
wire n_3175;
wire n_4594;
wire n_3130;
wire n_3231;
wire n_4800;
wire n_1417;
wire n_4799;
wire n_5054;
wire u6_mem_b1_b_88;
wire n_5112;
wire n_2697;
wire n_5057;
wire n_5145;
wire n_3242;
wire n_4388;
wire u8_mem_b1_b_71;
wire n_4387;
wire n_2028;
wire n_4796;
wire n_1424;
wire n_4795;
wire n_5056;
wire u6_mem_b3_b_146;
wire n_5100;
wire n_3180;
wire n_4589;
wire n_3215;
wire n_3214;
wire n_4590;
wire n_3536;
wire n_2312;
wire n_5527;
wire n_5526;
wire n_4675;
wire n_5381;
wire u11_mem_b1_b_149;
wire n_5300;
wire n_6502;
wire n_5052;
wire u6_mem_b3_b_143;
wire n_3169;
wire n_5053;
wire u6_mem_b3_b_144;
wire n_3228;
wire n_10902;
wire n_10206;
wire n_7241;
wire n_7089;
wire n_12504;
wire n_10201;
wire n_12483;
wire n_7084;
wire n_10202;
wire n_7239;
wire n_7085;
wire n_12161;
wire n_10199;
wire n_7235;
wire n_7181;
wire n_10200;
wire n_7236;
wire n_7182;
wire n_10196;
wire n_7232;
wire n_7178;
wire n_10198;
wire n_7233;
wire n_7179;
wire n_11721;
wire u3_mem_b0_b_101;
wire n_6522;
wire u11_mem_b1_b;
wire o7_status;
wire n_5618;
wire u6_mem_b2_b_47;
wire n_9137;
wire n_3865;
wire n_2763;
wire u6_mem_b3_b_132;
wire n_9109;
wire n_5952;
wire n_5951;
wire n_5987;
wire u4_mem_b1_b_84;
wire n_8322;
wire n_10922;
wire n_552;
wire n_4402;
wire u8_mem_b1_b_62;
wire n_4502;
wire n_2058;
wire n_1285;
wire n_1262;
wire u11_mem_b3_b_80;
wire n_10852;
wire n_2055;
wire n_2054;
wire n_2732;
wire n_2053;
wire n_2684;
wire n_2118;
wire n_2056;
wire n_1985;
wire n_2728;
wire n_2788;
wire n_2748;
wire n_2731;
wire n_2784;
wire n_2730;
wire n_2751;
wire n_2804;
wire n_2057;
wire n_2734;
wire n_1226;
wire u6_mem_b0_b_111;
wire n_8768;
wire n_2727;
wire n_1147;
wire n_2765;
wire n_1632;
wire n_2477;
wire n_4001;
wire n_1567;
wire n_1566;
wire n_910;
wire u26_ps_cnt_b3_b;
wire n_760;
wire n_1120;
wire n_11762;
wire n_1119;
wire n_550;
wire u13_ints_r_b7_b;
wire n_488;
wire n_3955;
wire n_5371;
wire n_6393;
wire n_6392;
wire n_6856;
wire n_6391;
wire n_6390;
wire n_6586;
wire n_6389;
wire n_6388;
wire n_6453;
wire n_6017;
wire n_5960;
wire n_5959;
wire n_5997;
wire n_6387;
wire n_6386;
wire n_6602;
wire n_6385;
wire n_6384;
wire n_6599;
wire n_6383;
wire n_6382;
wire n_6596;
wire n_6381;
wire n_6380;
wire n_6592;
wire n_6378;
wire n_6377;
wire n_6521;
wire n_6271;
wire n_5707;
wire n_6318;
wire n_5905;
wire n_2567;
wire n_6275;
wire n_6159;
wire n_12046;
wire n_6204;
wire n_3472;
wire n_12369;
wire u6_mem_b0_b_118;
wire n_5831;
wire n_10940;
wire n_2343;
wire n_459;
wire oc0_cfg;
wire n_10794;
wire n_10341;
wire n_9968;
wire n_9620;
wire i4_full;
wire n_608;
wire n_1157;
wire n_487;
wire n_10904;
wire n_10795;
wire n_11105;
wire n_6773;
wire n_12503;
wire n_1481;
wire n_10796;
wire n_9534;
wire n_668;
wire n_10905;
wire n_10342;
wire n_9694;
wire i3_full;
wire n_9690;
wire n_739;
wire n_9758;
wire n_9532;
wire n_10483;
wire n_611;
wire n_10928;
wire n_12006;
wire n_12007;
wire n_1473;
wire n_10801;
wire n_9964;
wire n_11600;
wire n_5624;
wire n_5632;
wire n_1777;
wire n_1833;
wire n_6838;
wire n_814;
wire n_415;
wire u2_res_cnt_b1_b;
wire u2_res_cnt_b3_b;
wire n_10934;
wire n_12012;
wire n_12013;
wire n_10791;
wire n_10998;
wire n_10789;
wire n_10933;
wire n_12140;
wire n_11536;
wire n_10932;
wire n_12150;
wire n_11538;
wire n_10931;
wire n_12042;
wire n_12043;
wire n_10930;
wire n_11950;
wire n_11951;
wire n_10945;
wire n_10929;
wire n_11980;
wire n_11981;
wire n_1010;
wire n_620;
wire n_1009;
wire n_531;
wire u11_mem_b1_b_124;
wire n_3952;
wire n_12818;
wire n_1124;
wire u14_n_134;
wire n_1755;
wire u11_mem_b0_b_171;
wire n_1425;
wire n_1924;
wire wb_din_673;
wire u7_mem_b0_b_104;
wire n_9400;
wire n_1158;
wire n_1008;
wire n_539;
wire u5_mem_b0_b_116;
wire n_8793;
wire n_509;
wire u9_mem_b2_b;
wire n_6463;
wire u10_mem_b1_b_130;
wire u11_mem_b3_b_83;
wire n_6182;
wire n_11453;
wire n_11454;
wire n_3374;
wire n_2391;
wire n_4646;
wire n_5480;
wire n_3492;
wire n_1260;
wire n_843;
wire u6_mem_b2_b_35;
wire n_9115;
wire u4_mem_b3_b_125;
wire i3_dout_575;
wire n_4064;
wire u5_mem_b2_b_30;
wire n_9247;
wire u6_mem_b3_b_140;
wire n_9099;
wire u4_mem_b1_b_77;
wire n_8332;
wire u5_mem_b3_b_126;
wire n_9203;
wire n_5063;
wire u6_mem_b3_b_152;
wire n_3022;
wire u6_mem_b0_b_119;
wire n_8761;
wire n_2692;
wire n_2721;
wire n_920;
wire u3_mem_b1_b_76;
wire n_8888;
wire n_2001;
wire n_938;
wire n_2707;
wire u8_mem_b2_b_42;
wire n_8881;
wire n_473;
wire n_751;
wire n_3934;
wire u9_din_tmp_55;
wire n_2368;
wire n_3935;
wire n_1498;
wire n_2831;
wire n_1409;
wire n_3087;
wire u5_mem_b1_b_86;
wire n_2281;
wire u7_mem_b0_b_100;
wire n_2282;
wire u6_mem_b2_b_39;
wire n_2285;
wire i6_empty;
wire n_5383;
wire n_11708;
wire u6_mem_b1_b_70;
wire u7_mem_b1_b_81;
wire n_9046;
wire n_5591;
wire n_2284;
wire n_1999;
wire n_2470;
wire n_5107;
wire u4_mem_b3_b_131;
wire n_5106;
wire n_2882;
wire n_4165;
wire u6_mem_b1_b_83;
wire n_9383;
wire u8_mem_b0_b_102;
wire n_3817;
wire n_7490;
wire n_9385;
wire u8_mem_b0_b_101;
wire n_3814;
wire n_8720;
wire u3_mem_b0_b_107;
wire n_3815;
wire n_8700;
wire n_8721;
wire n_3602;
wire n_9386;
wire u8_mem_b0_b;
wire n_3604;
wire n_8722;
wire u3_mem_b0_b_106;
wire n_3603;
wire n_7423;
wire n_9387;
wire u3_mem_b0_b_105;
wire n_3804;
wire n_8252;
wire u3_mem_b0_b_104;
wire n_3813;
wire n_3933;
wire u9_din_tmp_56;
wire u6_mem_b0_b_97;
wire n_9404;
wire n_977;
wire n_8718;
wire u8_mem_b0_b_103;
wire n_3818;
wire n_8719;
wire n_3601;
wire u6_mem_b1_b_78;
wire n_9177;
wire n_8014;
wire u4_mem_b2_b_41;
wire n_9250;
wire n_4359;
wire n_9212;
wire n_7884;
wire n_8013;
wire u4_mem_b2_b_42;
wire n_5443;
wire n_4087;
wire n_8012;
wire u4_mem_b2_b_43;
wire u6_wp_b2_b;
wire n_9465;
wire n_8228;
wire n_6681;
wire n_7462;
wire u14_u3_full_empty_r;
wire n_9537;
wire u10_mem_b3_b_85;
wire n_10682;
wire n_4853;
wire n_2615;
wire u2_to_cnt_b5_b;
wire n_2616;
wire n_8010;
wire u4_mem_b2_b_45;
wire n_2977;
wire n_7299;
wire i4_dout_622;
wire n_5355;
wire n_3339;
wire n_4135;
wire n_2974;
wire n_11789;
wire u8_mem_b0_b_119;
wire n_8009;
wire u4_mem_b2_b_46;
wire n_2253;
wire u8_mem_b2_b_45;
wire n_2362;
wire n_7202;
wire n_5728;
wire n_6815;
wire n_3698;
wire u5_mem_b0_b_121;
wire n_3720;
wire n_2251;
wire u4_mem_b3_b_124;
wire n_3697;
wire wb_din_663;
wire n_8992;
wire n_4541;
wire n_7663;
wire n_8993;
wire n_4538;
wire n_7664;
wire n_8995;
wire n_4536;
wire n_8145;
wire n_8996;
wire n_4309;
wire n_7665;
wire n_8988;
wire n_4366;
wire n_8948;
wire n_7658;
wire n_8989;
wire n_4339;
wire n_7659;
wire n_8990;
wire n_4546;
wire n_7660;
wire n_8991;
wire n_4307;
wire n_8981;
wire n_7661;
wire n_7303;
wire n_6700;
wire n_7110;
wire n_8986;
wire n_4292;
wire n_7656;
wire n_8987;
wire n_4305;
wire n_7657;
wire n_7386;
wire i3_dout_588;
wire n_7106;
wire n_3707;
wire u5_mem_b0_b_118;
wire wb_din_688;
wire u8_mem_b1_b_90;
wire n_8351;
wire i4_dout_620;
wire n_7045;
wire n_3704;
wire u5_mem_b0_b_119;
wire n_841;
wire n_7300;
wire i4_dout_621;
wire n_7109;
wire n_3700;
wire u5_mem_b0_b_92;
wire wb_din_662;
wire u10_mem_b3_b_77;
wire n_10694;
wire n_6448;
wire u11_mem_b2_b_89;
wire n_3699;
wire u5_mem_b0_b_120;
wire n_4627;
wire n_2459;
wire n_2636;
wire n_6920;
wire n_4621;
wire n_3351;
wire n_3712;
wire u5_mem_b0_b_115;
wire n_3710;
wire u7_mem_b0_b;
wire wb_din;
wire n_3709;
wire wb_din_686;
wire n_4730;
wire n_4729;
wire oc4_cfg_1004;
wire ic0_cfg_1024;
wire n_1862;
wire n_5998;
wire n_4882;
wire u7_mem_b3_b_144;
wire n_4961;
wire n_3324;
wire n_4728;
wire n_5277;
wire crac_out_865;
wire n_6972;
wire n_4727;
wire n_5272;
wire u13_intm_r_b20_b;
wire u13_ints_r_b20_b;
wire n_4726;
wire n_7488;
wire n_5196;
wire n_4236;
wire n_3104;
wire i6_dout_627;
wire n_4009;
wire n_5119;
wire u7_mem_b1_b_61;
wire n_5118;
wire n_2783;
wire n_4302;
wire u8_mem_b1_b_66;
wire n_2046;
wire n_2034;
wire n_2032;
wire n_945;
wire n_2772;
wire n_2714;
wire n_2713;
wire n_2035;
wire n_2103;
wire n_2744;
wire n_2036;
wire n_2792;
wire n_933;
wire u13_intm_r_b17_b;
wire u13_ints_r_b17_b;
wire n_2039;
wire n_2767;
wire n_2037;
wire n_2081;
wire n_4886;
wire u7_mem_b3_b_135;
wire n_2930;
wire n_1239;
wire n_1238;
wire n_5352;
wire n_2711;
wire u4_mem_b0_b_118;
wire n_8820;
wire u6_mem_b0_b_98;
wire n_8754;
wire n_2855;
wire u6_mem_b0_b_93;
wire u13_ints_r_b18_b;
wire n_6672;
wire u9_mem_b0_b_161;
wire n_10172;
wire n_8025;
wire u4_mem_b1_b_62;
wire n_2854;
wire n_2443;
wire u5_mem_b3_b_147;
wire n_12681;
wire n_12674;
wire n_12675;
wire n_12676;
wire n_12680;
wire n_2229;
wire u6_mem_b2_b;
wire u5_mem_b2_b_46;
wire n_11091;
wire n_12679;
wire u5_mem_b0_b_108;
wire n_12678;
wire n_12677;
wire n_1555;
wire n_1710;
wire n_6902;
wire n_6912;
wire n_11459;
wire u6_mem_b2_b_44;
wire n_9141;
wire n_2647;
wire n_1930;
wire n_2794;
wire n_2045;
wire n_1931;
wire n_2648;
wire n_1016;
wire n_1934;
wire n_2085;
wire n_1935;
wire n_2006;
wire n_1932;
wire n_2171;
wire n_2818;
wire n_1933;
wire n_5150;
wire u3_mem_b1_b_66;
wire n_5157;
wire n_2651;
wire n_5149;
wire n_2781;
wire n_3889;
wire u8_mem_b3_b_134;
wire n_1458;
wire n_5154;
wire u3_mem_b1_b_62;
wire n_2789;
wire n_5153;
wire u3_mem_b1_b_63;
wire n_2718;
wire u7_mem_b2_b_58;
wire n_4540;
wire n_2222;
wire n_5152;
wire u3_mem_b1_b_64;
wire n_2679;
wire n_4539;
wire u6_mem_b2_b_52;
wire n_4544;
wire n_2219;
wire n_5151;
wire u3_mem_b1_b_65;
wire n_2776;
wire n_3888;
wire u8_mem_b3_b_141;
wire n_1504;
wire n_4593;
wire n_3528;
wire n_2235;
wire n_10914;
wire n_11912;
wire n_12535;
wire u7_mem_b3_b_145;
wire n_8963;
wire u9_mem_b2_b_99;
wire n_10285;
wire u11_mem_b3_b_77;
wire n_10855;
wire n_10948;
wire n_10340;
wire n_11772;
wire n_2543;
wire n_196;
wire n_2542;
wire n_9092;
wire u4_mem_b0_b_111;
wire n_8825;
wire n_1706;
wire n_6893;
wire n_6905;
wire u2_to_cnt_b3_b;
wire n_6065;
wire n_1836;
wire n_6884;
wire n_6873;
wire u10_mem_b1_b_148;
wire n_10664;
wire n_5714;
wire n_5713;
wire u11_mem_b3_b_85;
wire n_10847;
wire n_5627;
wire u4_rp_b0_b;
wire n_10807;
wire n_2353;
wire u8_mem_b2_b_38;
wire n_6819;
wire n_6814;
wire n_9086;
wire n_5006;
wire n_9087;
wire n_7739;
wire n_9085;
wire n_5061;
wire n_7738;
wire n_6304;
wire n_6167;
wire n_6316;
wire n_5917;
wire n_5837;
wire n_5918;
wire n_5841;
wire n_5919;
wire n_9094;
wire n_9165;
wire n_7745;
wire n_9093;
wire n_7744;
wire n_9097;
wire n_5051;
wire n_7747;
wire n_9096;
wire n_4921;
wire n_7746;
wire n_9089;
wire n_4920;
wire n_7741;
wire n_8030;
wire u4_mem_b1_b_87;
wire n_9105;
wire n_7743;
wire n_9091;
wire n_7742;
wire n_10428;
wire n_5659;
wire n_1581;
wire n_10426;
wire n_5646;
wire n_10128;
wire n_5647;
wire n_1685;
wire n_10429;
wire n_5648;
wire n_1585;
wire n_10423;
wire n_5471;
wire n_10811;
wire n_9902;
wire n_10425;
wire n_10422;
wire n_10421;
wire n_5470;
wire n_1240;
wire u10_mem_b3_b_70;
wire n_10228;
wire n_12852;
wire n_3548;
wire n_3399;
wire n_5191;
wire n_3499;
wire n_3482;
wire n_4680;
wire n_3943;
wire n_5250;
wire n_4634;
wire n_5468;
wire u9_mem_b0_b_171;
wire n_4639;
wire n_5193;
wire n_3354;
wire n_2957;
wire n_5641;
wire n_5228;
wire n_5639;
wire u10_mem_b0_b_178;
wire n_5229;
wire u3_mem_b2_b_30;
wire n_8400;
wire n_2437;
wire n_3331;
wire n_4553;
wire n_2389;
wire n_2367;
wire n_1269;
wire n_763;
wire n_1790;
wire n_765;
wire n_1149;
wire n_1045;
wire n_969;
wire n_689;
wire u9_wp_b2_b;
wire u4_mem_b3_b_130;
wire n_9319;
wire n_1411;
wire oc1_cfg_976;
wire n_8569;
wire u11_din_tmp1;
wire n_10115;
wire n_6491;
wire n_6490;
wire n_5312;
wire n_6475;
wire n_6478;
wire n_6472;
wire n_6471;
wire n_6514;
wire n_5409;
wire n_6473;
wire n_2968;
wire n_3900;
wire u11_din_tmp_55;
wire n_4097;
wire oc3_int_set;
wire n_10091;
wire n_1203;
wire n_9951;
wire u10_mem_b2_b_109;
wire n_10768;
wire n_3899;
wire u10_din_tmp_55;
wire n_3911;
wire u6_mem_b1_b_73;
wire n_9187;
wire i3_status_1022;
wire n_5449;
wire n_5253;
wire u13_intm_r_b15_b;
wire crac_din_706;
wire n_4991;
wire u7_mem_b1_b_79;
wire u4_mem_b0_b_105;
wire n_8833;
wire n_6063;
wire n_1295;
wire n_6342;
wire n_6578;
wire n_5374;
wire u9_mem_b3_b_77;
wire n_925;
wire oc0_cfg_966;
wire n_7625;
wire u7_mem_b3_b_125;
wire n_7651;
wire n_7624;
wire u7_mem_b3_b_126;
wire u10_mem_b0_b_162;
wire n_7629;
wire u8_mem_b3_b_137;
wire n_7628;
wire u7_mem_b3_b_151;
wire n_7627;
wire u7_mem_b3_b_152;
wire n_7626;
wire u7_mem_b3_b_124;
wire n_7633;
wire u7_mem_b3_b_148;
wire n_7632;
wire u7_mem_b3_b_149;
wire n_7631;
wire u7_mem_b3_b_150;
wire n_7630;
wire u7_mem_b3_b_123;
wire u14_u7_full_empty_r;
wire n_7557;
wire n_9796;
wire n_8190;
wire n_8191;
wire o7_we;
wire n_7020;
wire n_9352;
wire in_valid_s_b0_b;
wire n_1308;
wire n_8660;
wire n_12585;
wire n_7537;
wire n_12335;
wire n_8661;
wire n_9475;
wire n_8662;
wire n_5825;
wire n_7538;
wire n_8663;
wire n_5382;
wire n_2563;
wire n_3930;
wire n_1593;
wire n_1590;
wire u4_mem_b2_b_48;
wire n_8287;
wire n_4015;
wire n_1616;
wire n_1613;
wire n_4014;
wire n_1611;
wire n_1607;
wire n_4808;
wire n_2525;
wire n_2523;
wire n_4013;
wire n_1606;
wire n_1603;
wire n_4012;
wire n_1601;
wire n_1855;
wire n_5705;
wire n_6161;
wire n_2927;
wire n_2924;
wire n_3143;
wire n_2402;
wire n_4011;
wire n_1597;
wire n_1594;
wire n_2516;
wire u10_mem_b2_b_116;
wire n_10752;
wire u11_mem_b2_b_113;
wire n_10866;
wire n_4995;
wire u5_mem_b3_b_135;
wire n_2934;
wire u9_mem_b3_b_76;
wire n_10711;
wire n_2519;
wire n_2344;
wire ac97_reset_pad_o_;
wire n_9491;
wire u4_mem_b3_b_132;
wire n_8262;
wire n_12588;
wire n_4829;
wire n_2568;
wire u9_rp_b0_b;
wire n_7369;
wire valid_s;
wire n_12590;
wire n_10663;
wire n_12340;
wire n_12336;
wire n_12592;
wire n_11128;
wire n_12591;
wire n_12370;
wire n_12368;
wire n_12361;
wire n_12362;
wire n_12363;
wire n_12367;
wire n_11846;
wire u4_mem_b3_b_136;
wire n_12744;
wire n_12273;
wire u4_mem_b1_b_74;
wire n_10742;
wire n_6866;
wire u9_mem_b0_b_165;
wire n_2517;
wire n_7581;
wire u3_mem_b1_b_77;
wire u4_mem_b3_b_140;
wire n_9345;
wire u4_mem_b1_b_89;
wire n_8313;
wire n_8454;
wire n_3847;
wire n_8452;
wire n_8097;
wire n_8158;
wire n_8462;
wire n_3842;
wire n_8460;
wire n_8911;
wire n_8164;
wire n_8032;
wire u4_mem_b1_b_85;
wire n_8463;
wire n_5155;
wire n_8026;
wire u4_mem_b1_b_90;
wire n_8230;
wire n_6684;
wire n_7464;
wire n_8459;
wire n_8163;
wire n_8027;
wire n_10743;
wire n_8446;
wire u7_mem_b2_b_41;
wire n_4509;
wire n_1995;
wire u7_mem_b2_b_39;
wire n_2064;
wire n_4890;
wire u7_mem_b1_b_68;
wire n_2688;
wire n_4319;
wire u8_mem_b1_b_87;
wire n_1946;
wire n_11029;
wire u3_mem_b3_b_133;
wire n_5133;
wire n_2912;
wire u7_mem_b2_b_42;
wire n_2060;
wire n_4312;
wire u7_mem_b2_b_53;
wire n_4313;
wire u7_mem_b2_b_47;
wire n_1944;
wire n_4441;
wire u4_mem_b2_b_38;
wire n_4439;
wire n_1947;
wire n_8613;
wire n_4687;
wire n_8611;
wire u7_mem_b1_b_72;
wire n_9061;
wire n_12371;
wire n_12066;
wire n_12111;
wire n_3317;
wire n_2914;
wire n_3396;
wire n_2467;
wire u5_mem_b1_b_61;
wire n_9287;
wire n_4586;
wire n_3537;
wire n_2897;
wire n_5032;
wire u5_mem_b1_b_79;
wire n_5037;
wire n_2778;
wire n_10613;
wire n_6265;
wire n_6229;
wire n_10617;
wire n_5033;
wire u5_mem_b1_b_60;
wire n_2661;
wire n_5034;
wire u5_mem_b1_b_78;
wire n_2799;
wire n_5035;
wire u5_mem_b1_b_77;
wire n_2666;
wire n_5036;
wire u6_mem_b3_b_137;
wire n_3296;
wire n_5038;
wire u5_mem_b1_b_76;
wire n_2726;
wire n_5039;
wire u5_mem_b1_b_75;
wire n_5048;
wire n_2779;
wire n_5040;
wire u5_mem_b1_b_74;
wire n_2747;
wire n_5041;
wire u6_mem_b3_b_138;
wire n_3357;
wire n_11619;
wire n_7123;
wire n_7069;
wire n_11617;
wire n_7216;
wire n_6983;
wire n_10496;
wire n_7219;
wire n_7067;
wire n_10481;
wire n_11615;
wire n_7121;
wire n_7064;
wire n_10493;
wire n_7217;
wire n_7066;
wire n_11633;
wire n_7218;
wire n_6984;
wire n_7476;
wire n_6745;
wire n_7337;
wire n_7383;
wire n_6718;
wire n_11564;
wire n_11534;
wire n_1230;
wire n_7030;
wire n_7365;
wire n_7050;
wire n_5965;
wire n_2271;
wire n_4306;
wire u5_mem_b2_b_32;
wire n_4370;
wire n_2134;
wire u11_mem_b1_b_123;
wire n_10549;
wire n_7450;
wire n_6692;
wire n_7302;
wire crac_out_864;
wire n_8631;
wire n_7479;
wire in_valid_s_b1_b;
wire n_4247;
wire u7_mem_b1_b_75;
wire n_7478;
wire n_7477;
wire i3_dout_568;
wire n_4042;
wire oc1_cfg_979;
wire n_8564;
wire out_slt_65;
wire n_11101;
wire n_4442;
wire u4_mem_b2_b;
wire n_2106;
wire n_2638;
wire u8_mem_b2_b_51;
wire n_3441;
wire n_3224;
wire u5_mem_b0_b_117;
wire n_3225;
wire n_12840;
wire u4_mem_b0_b_113;
wire u8_mem_b2_b_52;
wire n_4491;
wire n_1826;
wire n_4333;
wire n_214;
wire u9_din_tmp_49;
wire n_9771;
wire n_5494;
wire u11_mem_b3_b_76;
wire u9_mem_b0_b_157;
wire n_10142;
wire n_10108;
wire n_4443;
wire n_2023;
wire n_5890;
wire n_5823;
wire n_6152;
wire n_6397;
wire n_6396;
wire n_6582;
wire n_6867;
wire n_6883;
wire n_4927;
wire u6_mem_b3_b_131;
wire n_2916;
wire n_12531;
wire n_6869;
wire n_6868;
wire n_6925;
wire n_6812;
wire n_6407;
wire n_6406;
wire n_6563;
wire n_6401;
wire n_6400;
wire n_6539;
wire n_6399;
wire n_6398;
wire n_6405;
wire n_6404;
wire n_6646;
wire n_6810;
wire n_6797;
wire n_3515;
wire n_12067;
wire n_12379;
wire oc3_cfg_996;
wire n_8542;
wire u9_din_tmp1;
wire n_9789;
wire n_5550;
wire n_12626;
wire n_670;
wire n_921;
wire n_481;
wire u10_rp_b1_b;
wire u10_rp_b0_b;
wire n_2369;
wire n_1111;
wire n_673;
wire n_980;
wire u13_ints_r_b0_b;
wire n_1036;
wire n_12281;
wire n_244;
wire u8_mem_b1_b_60;
wire n_8926;
wire u9_mem_b2_b_95;
wire n_10265;
wire n_672;
wire n_671;
wire n_924;
wire u11_mem_b0_b_158;
wire n_10413;
wire n_5563;
wire n_5884;
wire u10_din_tmp_42;
wire n_9853;
wire u7_mem_b2_b_46;
wire n_4232;
wire n_7373;
wire n_11037;
wire n_4525;
wire n_2211;
wire u7_mem_b2_b_56;
wire n_2878;
wire u3_mem_b2_b_34;
wire n_3207;
wire u10_din_tmp_50;
wire n_9862;
wire n_5877;
wire n_5879;
wire n_5876;
wire n_9103;
wire n_7752;
wire n_12195;
wire n_12196;
wire n_11069;
wire n_11060;
wire n_12064;
wire n_12065;
wire n_11059;
wire n_11145;
wire n_10982;
wire n_11144;
wire n_11062;
wire n_12193;
wire n_12194;
wire n_11056;
wire n_10607;
wire n_10188;
wire n_11055;
wire n_11743;
wire n_11744;
wire n_5839;
wire n_11058;
wire n_10609;
wire n_12505;
wire n_11057;
wire n_12793;
wire n_12794;
wire n_3124;
wire u7_mem_b1_b_66;
wire n_3522;
wire n_3125;
wire u6_mem_b0_b_108;
wire n_11054;
wire n_12543;
wire n_11746;
wire n_11053;
wire n_11749;
wire n_11750;
wire n_740;
wire n_6752;
wire n_6751;
wire n_495;
wire u9_mem_b3_b_85;
wire n_10702;
wire n_8705;
wire u8_mem_b0_b_111;
wire n_3831;
wire n_8707;
wire u8_mem_b0_b_110;
wire n_3830;
wire n_8703;
wire n_3836;
wire n_8704;
wire u8_mem_b0_b_112;
wire n_3833;
wire n_8699;
wire u8_mem_b0_b_114;
wire n_3838;
wire n_3592;
wire n_8696;
wire u3_mem_b0_b_114;
wire n_3627;
wire n_8698;
wire u8_mem_b0_b_115;
wire n_3590;
wire u7_mem_b2_b_43;
wire n_9379;
wire u8_mem_b0_b_116;
wire n_3589;
wire u9_mem_b2_b_90;
wire n_10272;
wire n_11041;
wire u11_mem_b1_b_125;
wire n_9330;
wire n_5078;
wire n_7960;
wire n_762;
wire n_782;
wire crac_din_703;
wire n_1193;
wire u3_mem_b3_b_136;
wire n_8381;
wire u9_mem_b0_b_169;
wire n_10164;
wire u3_mem_b0_b_93;
wire n_8684;
wire n_8962;
wire n_4881;
wire n_8961;
wire n_7635;
wire n_4898;
wire n_7636;
wire n_8967;
wire n_4883;
wire n_7639;
wire n_8968;
wire n_5159;
wire n_7640;
wire n_8964;
wire n_7637;
wire n_8965;
wire n_5073;
wire n_7638;
wire n_8972;
wire n_4952;
wire n_8971;
wire n_7643;
wire n_8973;
wire n_5076;
wire n_7644;
wire n_8969;
wire n_4884;
wire n_7641;
wire n_8970;
wire n_7642;
wire n_4529;
wire n_1948;
wire n_2127;
wire n_2120;
wire n_2829;
wire u6_mem_b0_b_101;
wire n_8779;
wire n_4528;
wire u3_mem_b2_b_43;
wire n_4533;
wire n_2079;
wire n_2130;
wire n_2083;
wire n_2782;
wire n_1499;
wire n_4489;
wire u8_mem_b2_b_33;
wire n_1805;
wire u11_mem_b1_b_137;
wire n_10896;
wire u3_mem_b2_b_41;
wire n_8421;
wire dma_req_o_b3_b;
wire n_11193;
wire n_10839;
wire n_9905;
wire n_10391;
wire n_9818;
wire n_9721;
wire n_9674;
wire n_2021;
wire n_2020;
wire n_2704;
wire n_2775;
wire n_3878;
wire u8_mem_b3_b_143;
wire n_1479;
wire n_2701;
wire u10_mem_b1_b_144;
wire n_10805;
wire n_4377;
wire u5_mem_b2_b_38;
wire n_4378;
wire n_2699;
wire n_1827;
wire n_2698;
wire n_2716;
wire n_2018;
wire n_3350;
wire u9_mem_b2_b_110;
wire n_10725;
wire n_888;
wire n_4488;
wire u6_mem_b2_b_41;
wire n_4504;
wire n_1952;
wire n_3347;
wire n_11963;
wire n_10645;
wire n_11977;
wire n_2657;
wire n_2761;
wire n_1943;
wire n_2735;
wire n_2658;
wire n_6670;
wire n_461;
wire n_6510;
wire n_3717;
wire u5_mem_b0_b_112;
wire wb_din_682;
wire n_1495;
wire n_11959;
wire n_11997;
wire n_11961;
wire n_4836;
wire n_1404;
wire n_9777;
wire n_9642;
wire n_2653;
wire n_9514;
wire n_4500;
wire n_4499;
wire n_2004;
wire n_4498;
wire u6_mem_b2_b_43;
wire n_1984;
wire n_4501;
wire u7_mem_b2_b_48;
wire n_1964;
wire u13_intm_r_b2_b;
wire n_8494;
wire n_3884;
wire u8_mem_b3_b_136;
wire n_1423;
wire u8_mem_b3_b_135;
wire n_8458;
wire n_5128;
wire u7_mem_b1_b_77;
wire n_2722;
wire n_5127;
wire u3_mem_b3_b_123;
wire n_3067;
wire n_4496;
wire u7_mem_b2_b_29;
wire n_5126;
wire u3_mem_b3_b_130;
wire n_3512;
wire u9_mem_b0_b_177;
wire n_10155;
wire u26_ps_cnt_b5_b;
wire n_9593;
wire n_2578;
wire u13_ints_r_b15_b;
wire n_3985;
wire u9_mem_b3_b_70;
wire n_10256;
wire u16_u8_dma_req_r1;
wire n_11907;
wire n_2953;
wire n_9469;
wire ic2_int_set;
wire n_9545;
wire n_2506;
wire u7_mem_b3_b_133;
wire n_8979;
wire n_3674;
wire wb_din_678;
wire n_3671;
wire u6_mem_b0_b_113;
wire n_3676;
wire u6_mem_b0_b_105;
wire wb_din_675;
wire n_3675;
wire u6_mem_b0_b_106;
wire wb_din_676;
wire n_3679;
wire u6_mem_b0_b_103;
wire n_3677;
wire wb_din_670;
wire n_3682;
wire u6_mem_b0_b_100;
wire n_813;
wire n_3681;
wire u6_mem_b0_b_102;
wire n_3670;
wire u6_mem_b0_b_116;
wire n_1060;
wire n_851;
wire i6_dout_649;
wire n_3826;
wire n_58;
wire n_178;
wire n_2625;
wire n_2624;
wire n_2621;
wire n_4081;
wire n_1291;
wire n_5941;
wire n_6326;
wire n_6266;
wire n_8205;
wire n_5588;
wire n_802;
wire n_806;
wire n_544;
wire oc2_cfg_986;
wire n_712;
wire n_145;
wire u4_rp_b3_b;
wire n_650;
wire n_10440;
wire n_5666;
wire n_1615;
wire n_9502;
wire n_7164;
wire n_9500;
wire n_7163;
wire n_10444;
wire n_5664;
wire n_1628;
wire n_10443;
wire n_5655;
wire n_9506;
wire n_7166;
wire n_1122;
wire n_12847;
wire n_9563;
wire n_7289;
wire n_1127;
wire n_12845;
wire n_9994;
wire n_1700;
wire n_10054;
wire n_9842;
wire n_5772;
wire n_9996;
wire n_10327;
wire n_771;
wire u4_mem_b2_b_44;
wire n_8294;
wire n_12801;
wire n_5656;
wire n_1072;
wire n_677;
wire u13_ints_r_b12_b;
wire n_676;
wire n_617;
wire u13_ints_r_b3_b;
wire n_616;
wire n_1384;
wire n_1605;
wire u11_mem_b0_b_175;
wire n_12136;
wire n_6079;
wire n_12532;
wire n_9292;
wire n_1701;
wire u9_mem_b0_b_174;
wire n_10923;
wire n_356;
wire u9_mem_b1_b_138;
wire n_6021;
wire u10_mem_b2_b_95;
wire n_1584;
wire u11_mem_b1_b_148;
wire n_598;
wire n_8197;
wire n_1199;
wire n_832;
wire n_931;
wire i6_dout_636;
wire n_4030;
wire u4_mem_b3_b_142;
wire n_9342;
wire n_811;
wire ic2_cfg_1044;
wire n_209;
wire u14_u8_full_empty_r;
wire n_10158;
wire u6_rp_b2_b;
wire n_11179;
wire n_118;
wire n_324;
wire n_465;
wire n_53;
wire u9_rp_b1_b;
wire n_4845;
wire u9_wp_b3_b;
wire u5_wp_b0_b;
wire n_9517;
wire n_6051;
wire n_5249;
wire n_303;
wire n_6716;
wire n_4846;
wire n_1818;
wire u2_res_cnt_b2_b;
wire n_7145;
wire n_6711;
wire n_7146;
wire n_8243;
wire n_6705;
wire n_7473;
wire n_12625;
wire n_3289;
wire u3_mem_b2_b_35;
wire n_8241;
wire n_4844;
wire n_7329;
wire i4_dout_617;
wire n_7133;
wire n_4028;
wire n_1665;
wire n_1664;
wire n_8242;
wire n_6677;
wire n_7472;
wire n_4812;
wire n_2531;
wire n_1236;
wire n_4024;
wire n_1654;
wire n_1652;
wire n_4026;
wire n_1658;
wire n_4025;
wire n_1656;
wire n_1655;
wire u5_mem_b1_b_87;
wire n_9291;
wire n_8424;
wire n_4532;
wire n_8393;
wire n_8138;
wire n_3856;
wire n_8133;
wire n_8075;
wire u3_mem_b3_b_127;
wire n_3227;
wire u3_mem_b2_b_47;
wire n_12619;
wire u4_mem_b3_b_149;
wire n_8071;
wire u3_mem_b2_b;
wire n_8238;
wire n_6676;
wire n_7461;
wire u7_mem_b2_b_34;
wire n_7736;
wire u6_mem_b3_b_151;
wire n_7735;
wire u6_mem_b3_b_150;
wire n_7737;
wire u6_mem_b3_b_123;
wire n_7740;
wire u6_mem_b3_b_148;
wire u6_mem_b3_b_149;
wire n_5060;
wire n_3220;
wire u11_mem_b2_b_101;
wire n_10529;
wire n_4198;
wire u7_mem_b1_b_86;
wire n_4130;
wire n_8431;
wire n_3885;
wire n_8146;
wire n_8430;
wire n_4348;
wire n_8144;
wire n_8428;
wire n_3854;
wire n_8143;
wire n_8427;
wire n_4534;
wire n_8440;
wire n_8142;
wire n_8054;
wire u4_mem_b1_b_70;
wire n_8233;
wire n_6688;
wire n_7467;
wire n_8434;
wire n_3883;
wire n_8148;
wire n_8432;
wire n_4537;
wire n_2448;
wire n_8045;
wire u4_mem_b1_b_76;
wire n_8044;
wire n_7988;
wire n_7987;
wire u4_mem_b2_b_37;
wire n_5302;
wire u9_mem_b3_b_81;
wire u8_mem_b0_b_109;
wire n_8709;
wire n_4901;
wire n_5069;
wire n_2674;
wire n_4902;
wire u7_mem_b1_b;
wire n_2671;
wire n_1322;
wire n_4905;
wire u7_mem_b1_b_69;
wire n_4903;
wire u7_mem_b1_b_73;
wire n_4904;
wire u7_mem_b1_b_71;
wire n_4907;
wire u7_mem_b3_b_132;
wire n_3079;
wire n_3849;
wire n_1484;
wire n_1485;
wire n_4320;
wire u3_mem_b2_b_52;
wire n_2121;
wire n_4906;
wire u6_mem_b1_b_68;
wire n_2659;
wire n_4393;
wire u8_mem_b1_b_89;
wire n_2005;
wire n_10780;
wire n_2067;
wire n_1180;
wire n_3229;
wire n_3259;
wire u5_mem_b0_b_104;
wire n_2865;
wire n_2487;
wire n_507;
wire n_12805;
wire u5_mem_b1_b_73;
wire n_3257;
wire n_5084;
wire u4_mem_b3_b_147;
wire n_5102;
wire n_2928;
wire n_4400;
wire u8_mem_b1_b_84;
wire n_2156;
wire u4_mem_b3_b_148;
wire n_3246;
wire n_5083;
wire n_2673;
wire u3_mem_b3_b_125;
wire n_8359;
wire n_2958;
wire u4_mem_b3_b_123;
wire n_2877;
wire u9_mem_b3_b_75;
wire n_10712;
wire n_6668;
wire u10_mem_b2_b_98;
wire n_12152;
wire n_6769;
wire n_10574;
wire n_6160;
wire n_5804;
wire n_9873;
wire n_9685;
wire n_12153;
wire n_6264;
wire n_11736;
wire n_10605;
wire n_11626;
wire n_10583;
wire u9_mem_b3_b_64;
wire n_10238;
wire n_11630;
wire n_5575;
wire u10_mem_b3_b_75;
wire n_9641;
wire n_12662;
wire n_5202;
wire n_4120;
wire n_2970;
wire u10_mem_b2_b_93;
wire n_10649;
wire n_12026;
wire n_12027;
wire n_1568;
wire n_6540;
wire n_9263;
wire u10_mem_b2_b_91;
wire n_10274;
wire u7_mem_b0_b_96;
wire n_192;
wire u7_mem_b3_b_127;
wire n_1538;
wire n_11853;
wire u7_mem_b1_b_65;
wire n_9695;
wire n_804;
wire i6_status_1042;
wire n_5638;
wire u4_wp_b2_b;
wire n_9468;
wire n_6793;
wire n_11925;
wire n_6443;
wire n_6441;
wire n_6440;
wire n_6439;
wire n_11542;
wire n_6794;
wire n_5973;
wire n_501;
wire n_6011;
wire n_6871;
wire n_5971;
wire n_406;
wire n_6449;
wire n_932;
wire n_6245;
wire n_6244;
wire n_6259;
wire n_6435;
wire n_6434;
wire n_6432;
wire n_2278;
wire n_8207;
wire n_564;
wire n_7327;
wire n_6123;
wire u9_mem_b3_b_57;
wire n_10251;
wire oc5_cfg_1020;
wire n_8195;
wire n_1381;
wire n_6714;
wire n_10092;
wire n_9769;
wire n_9601;
wire n_9661;
wire n_854;
wire n_510;
wire n_458;
wire n_3516;
wire u4_mem_b0_b_116;
wire n_10401;
wire n_9647;
wire n_9838;
wire n_10090;
wire n_9591;
wire n_9756;
wire n_7326;
wire n_6834;
wire n_6127;
wire n_12621;
wire n_12620;
wire n_5225;
wire n_593;
wire n_3159;
wire n_12825;
wire n_10088;
wire n_9587;
wire n_1791;
wire u5_mem_b2_b_48;
wire n_5586;
wire n_3976;
wire n_706;
wire n_1704;
wire u9_mem_b0_b_175;
wire n_10269;
wire n_6903;
wire n_10235;
wire i6_dout_656;
wire n_4007;
wire n_3162;
wire u6_mem_b0_b_112;
wire n_6864;
wire u9_mem_b0_b_166;
wire n_2507;
wire u9_mem_b0_b_179;
wire n_1786;
wire n_8188;
wire n_98;
wire u10_mem_b2_b_107;
wire n_11657;
wire u4_mem_b1_b_71;
wire n_12250;
wire n_6375;
wire u10_mem_b0_b_163;
wire n_3164;
wire n_5144;
wire u3_mem_b1_b_71;
wire n_2830;
wire n_2297;
wire u5_mem_b2_b_49;
wire n_3163;
wire n_3453;
wire n_4527;
wire n_2351;
wire n_5146;
wire u7_mem_b3_b_129;
wire n_3065;
wire n_913;
wire n_746;
wire n_705;
wire n_1108;
wire n_3106;
wire u7_mem_b2_b_33;
wire n_9490;
wire n_1887;
wire n_7533;
wire n_10623;
wire n_12144;
wire n_11077;
wire n_11962;
wire n_11976;
wire n_11075;
wire n_10626;
wire n_10209;
wire n_11081;
wire n_11956;
wire n_11957;
wire n_11083;
wire n_11080;
wire n_11958;
wire n_11079;
wire n_11996;
wire n_11078;
wire n_11960;
wire n_4390;
wire n_2062;
wire n_9368;
wire u3_mem_b0_b_95;
wire n_3771;
wire n_8682;
wire n_249;
wire u10_mem_b1_b_139;
wire n_1614;
wire u11_mem_b1_b_142;
wire n_5377;
wire u10_mem_b2_b_112;
wire n_8687;
wire u8_mem_b0_b_98;
wire n_3649;
wire n_8688;
wire u8_mem_b0_b_97;
wire n_3570;
wire n_8689;
wire u8_mem_b0_b_96;
wire n_3750;
wire n_9369;
wire u3_mem_b0_b_119;
wire n_3582;
wire n_3744;
wire n_8250;
wire n_8685;
wire u3_mem_b0_b_120;
wire n_3579;
wire n_8686;
wire u8_mem_b0_b_99;
wire n_3580;
wire n_4391;
wire n_1988;
wire i4_dout_625;
wire n_3998;
wire n_4596;
wire n_3240;
wire n_3238;
wire n_8934;
wire n_4392;
wire u3_mem_b2_b_58;
wire n_4519;
wire n_2086;
wire n_2952;
wire n_3252;
wire n_3486;
wire n_8984;
wire n_2954;
wire n_2955;
wire n_3423;
wire n_4597;
wire n_3176;
wire n_3071;
wire n_2331;
wire u7_mem_b0_b_105;
wire n_4125;
wire u7_mem_b1_b_74;
wire n_5379;
wire n_5290;
wire n_5424;
wire n_9000;
wire n_2951;
wire n_2200;
wire u7_mem_b0_b_106;
wire n_4828;
wire n_2610;
wire n_2587;
wire n_6140;
wire n_5709;
wire n_6091;
wire n_6143;
wire n_6142;
wire n_6141;
wire u10_mem_b0_b_156;
wire n_10120;
wire n_6139;
wire n_4629;
wire n_5200;
wire n_2619;
wire n_4633;
wire u11_mem_b1_b_147;
wire n_10882;
wire n_1172;
wire u3_wp_b1_b;
wire n_937;
wire n_8648;
wire n_1129;
wire n_2137;
wire n_10003;
wire n_5357;
wire n_10010;
wire n_2911;
wire u3_mem_b1_b_85;
wire n_3316;
wire n_9007;
wire n_11905;
wire dma_req_o_b8_b;
wire n_11903;
wire u16_u4_dma_req_r1;
wire n_11123;
wire n_2026;
wire n_2025;
wire u5_mem_b0_b_105;
wire n_8804;
wire n_9820;
wire n_2003;
wire n_2010;
wire n_2096;
wire n_2476;
wire n_867;
wire n_2012;
wire n_2099;
wire n_2011;
wire n_2041;
wire n_2007;
wire n_2009;
wire n_2008;
wire n_2693;
wire n_11904;
wire n_12743;
wire n_12742;
wire n_521;
wire u4_rp_b2_b;
wire n_12747;
wire n_12738;
wire n_602;
wire n_12739;
wire n_12740;
wire n_12741;
wire n_12745;
wire u4_mem_b0_b_103;
wire u4_mem_b3_b_134;
wire n_12755;
wire n_12748;
wire n_12749;
wire n_12750;
wire n_12754;
wire n_1449;
wire n_2662;
wire n_2773;
wire n_1959;
wire n_2189;
wire n_1958;
wire n_821;
wire n_2660;
wire n_1956;
wire n_1957;
wire n_1954;
wire n_2133;
wire n_1955;
wire u10_mem_b1_b_132;
wire n_10205;
wire n_4508;
wire n_4507;
wire n_2146;
wire u3_mem_b3_b_134;
wire n_2985;
wire n_4512;
wire n_1941;
wire n_4511;
wire u3_mem_b2_b_37;
wire n_2027;
wire u8_mem_b3_b_148;
wire n_1476;
wire n_4510;
wire u7_mem_b2_b_49;
wire n_1945;
wire n_4515;
wire u6_mem_b2_b_46;
wire n_2234;
wire n_4514;
wire u4_mem_b1_b_88;
wire n_5140;
wire n_2762;
wire n_4513;
wire n_2141;
wire u3_mem_b2_b_51;
wire n_8346;
wire u4_mem_b2_b_34;
wire n_8269;
wire u10_mem_b3_b_86;
wire n_10681;
wire n_9039;
wire n_5005;
wire n_7696;
wire u10_mem_b0_b_174;
wire u11_mem_b1_b_138;
wire n_10895;
wire n_4565;
wire n_2252;
wire n_4563;
wire n_4561;
wire n_2248;
wire n_3894;
wire n_3020;
wire n_5643;
wire u10_mem_b0_b_179;
wire n_5227;
wire n_6573;
wire n_4557;
wire n_2240;
wire n_1730;
wire n_365;
wire n_5369;
wire n_6570;
wire n_3928;
wire n_2305;
wire n_6566;
wire n_4550;
wire n_2334;
wire n_1731;
wire n_45;
wire n_1736;
wire n_198;
wire n_5343;
wire n_3063;
wire u3_mem_b0_b_103;
wire n_8724;
wire n_1739;
wire n_1738;
wire n_1737;
wire n_1745;
wire n_1744;
wire n_1743;
wire n_1742;
wire n_5294;
wire u3_mem_b1_b_89;
wire n_8408;
wire n_476;
wire n_9134;
wire n_9133;
wire n_4531;
wire n_4523;
wire n_7782;
wire n_9136;
wire n_4335;
wire n_9170;
wire n_7781;
wire n_9140;
wire n_4505;
wire n_9139;
wire n_7784;
wire n_9138;
wire n_9182;
wire n_7783;
wire n_9142;
wire n_7786;
wire n_4336;
wire n_7785;
wire n_9144;
wire n_7788;
wire n_9143;
wire n_4337;
wire n_7787;
wire u4_mem_b0_b_97;
wire n_9432;
wire n_6315;
wire n_6239;
wire n_5937;
wire n_5857;
wire n_6826;
wire n_6322;
wire n_6254;
wire n_6323;
wire n_12530;
wire n_11541;
wire n_6800;
wire n_6317;
wire n_6194;
wire n_6319;
wire n_6320;
wire n_5719;
wire n_6321;
wire n_6246;
wire n_10386;
wire n_1754;
wire n_10384;
wire n_1619;
wire n_995;
wire n_520;
wire n_9654;
wire n_9496;
wire n_9483;
wire n_9651;
wire n_9495;
wire n_9481;
wire n_9494;
wire n_5615;
wire ac97_rst_force;
wire n_9597;
wire n_10390;
wire n_1650;
wire n_10389;
wire n_1644;
wire n_10388;
wire n_1633;
wire n_10387;
wire n_339;
wire n_2613;
wire n_4718;
wire dma_req_o_b6_b;
wire n_12373;
wire n_3973;
wire crac_out_861;
wire n_2582;
wire u13_ints_r_b4_b;
wire n_5451;
wire n_1386;
wire n_4148;
wire n_5165;
wire n_2380;
wire n_3052;
wire n_5164;
wire n_3191;
wire n_3030;
wire n_5163;
wire n_3282;
wire n_3473;
wire n_3975;
wire u13_ints_r_b2_b;
wire n_3979;
wire n_5162;
wire n_3107;
wire n_2903;
wire u10_din_tmp_47;
wire u13_ints_r_b28_b;
wire n_9453;
wire n_5620;
wire n_9943;
wire n_12149;
wire n_12688;
wire n_2586;
wire n_4719;
wire n_5285;
wire u10_mem_b1_b_147;
wire n_5284;
wire n_9719;
wire n_319;
wire n_471;
wire i3_dout_585;
wire n_4053;
wire n_6025;
wire n_5404;
wire u5_mem_b3_b_148;
wire n_9213;
wire n_6894;
wire n_6168;
wire n_12115;
wire n_6169;
wire n_6155;
wire n_5810;
wire n_5809;
wire n_5976;
wire n_5403;
wire n_6173;
wire n_6172;
wire n_11986;
wire n_6174;
wire n_6177;
wire n_6176;
wire n_12664;
wire n_6179;
wire n_11898;
wire n_6181;
wire n_6180;
wire n_4204;
wire u7_mem_b1_b_62;
wire n_9306;
wire u11_mem_b2_b_99;
wire u10_mem_b3_b_84;
wire n_6561;
wire n_6560;
wire n_6559;
wire u11_mem_b0_b_152;
wire n_6466;
wire n_4182;
wire u6_mem_b1_b_81;
wire u3_mem_b2_b_36;
wire n_3142;
wire u6_mem_b0_b_92;
wire n_11464;
wire u8_mem_b1_b_63;
wire n_12295;
wire n_3144;
wire u8_mem_b2_b_59;
wire u7_mem_b0_b_102;
wire n_11514;
wire u6_mem_b1_b_61;
wire n_10714;
wire n_4768;
wire n_10738;
wire n_10030;
wire n_10715;
wire n_4765;
wire n_10019;
wire n_10031;
wire n_4758;
wire n_10040;
wire n_10727;
wire n_10747;
wire n_10041;
wire n_10722;
wire n_4756;
wire n_10723;
wire n_4775;
wire n_10038;
wire n_10719;
wire n_4744;
wire n_10035;
wire n_10721;
wire n_4774;
wire n_10037;
wire n_10717;
wire n_4770;
wire n_10032;
wire n_10718;
wire n_4773;
wire n_10034;
wire n_4094;
wire u2_res_cnt_b0_b;
wire n_10074;
wire n_174;
wire n_10073;
wire n_10072;
wire n_9;
wire n_10065;
wire n_10076;
wire n_366;
wire n_10075;
wire n_349;
wire n_10068;
wire n_12339;
wire n_1096;
wire n_10067;
wire n_10071;
wire n_10069;
wire n_10066;
wire n_2545;
wire n_10064;
wire n_204;
wire n_10045;
wire n_11587;
wire n_11579;
wire n_11586;
wire u6_rp_b1_b;
wire u3_mem_b1_b_61;
wire n_8471;
wire n_7460;
wire i4_dout_608;
wire n_7297;
wire n_7348;
wire i4_dout_607;
wire n_7349;
wire i4_dout_603;
wire n_7340;
wire n_7149;
wire i4_dout_604;
wire n_7339;
wire u9_mem_b0_b_180;
wire n_10150;
wire n_7031;
wire i4_status;
wire i4_status_1032;
wire n_12828;
wire n_2777;
wire n_7280;
wire n_7018;
wire n_7363;
wire n_7148;
wire ic1_int_set_721;
wire n_5863;
wire n_11441;
wire n_3202;
wire n_11442;
wire n_4031;
wire n_1837;
wire n_1653;
wire n_11148;
wire n_5710;
wire n_2243;
wire n_3206;
wire n_3205;
wire n_2439;
wire n_5558;
wire n_5711;
wire n_6241;
wire n_11966;
wire n_3218;
wire n_11967;
wire n_2406;
wire n_5874;
wire n_12857;
wire n_12858;
wire n_11482;
wire n_1336;
wire n_5559;
wire n_3542;
wire n_3212;
wire n_2857;
wire n_2231;
wire oc3_cfg_997;
wire n_8540;
wire n_4606;
wire n_3551;
wire n_3297;
wire u4_mem_b1_b_73;
wire n_8340;
wire u5_mem_b2_b_40;
wire n_9270;
wire n_10946;
wire n_8801;
wire u11_mem_b3_b_60;
wire n_10452;
wire n_8835;
wire u4_mem_b0_b_102;
wire n_3799;
wire n_7499;
wire n_9442;
wire n_3797;
wire n_9441;
wire u4_mem_b0_b_104;
wire n_3796;
wire n_3795;
wire n_9443;
wire n_3811;
wire n_8838;
wire u4_mem_b0_b_100;
wire n_3802;
wire n_8837;
wire u4_mem_b0_b;
wire n_3803;
wire n_8836;
wire u4_mem_b0_b_101;
wire n_3801;
wire n_9440;
wire u4_mem_b0_b_106;
wire n_3791;
wire n_8832;
wire u4_mem_b0_b_107;
wire n_3788;
wire n_798;
wire n_710;
wire n_8949;
wire n_8005;
wire u4_mem_b2_b_49;
wire n_8004;
wire u4_mem_b2_b_50;
wire n_8003;
wire u4_mem_b2_b_51;
wire n_8002;
wire u4_mem_b2_b_52;
wire n_7287;
wire n_7443;
wire n_8643;
wire n_7518;
wire u4_mem_b0_b_120;
wire n_8816;
wire n_6678;
wire n_6686;
wire i6_dout_642;
wire i3_dout_580;
wire u6_mem_b2_b_57;
wire n_9124;
wire n_3318;
wire n_8405;
wire i6_dout_643;
wire i3_dout_581;
wire n_3684;
wire n_2329;
wire n_8839;
wire u3_mem_b0_b_109;
wire n_3823;
wire n_9035;
wire n_8841;
wire u3_mem_b0_b_118;
wire n_3584;
wire n_5103;
wire n_3307;
wire n_5104;
wire u4_mem_b3_b_133;
wire n_3309;
wire i6_dout_634;
wire i3_dout_572;
wire n_1039;
wire n_638;
wire n_4408;
wire n_1973;
wire n_5108;
wire n_2753;
wire n_4407;
wire n_2209;
wire out_slt_84;
wire n_10955;
wire n_8788;
wire n_4405;
wire n_1673;
wire n_5105;
wire n_3343;
wire n_8846;
wire n_5160;
wire n_8068;
wire n_6554;
wire u11_mem_b3_b;
wire n_707;
wire n_7771;
wire n_7768;
wire u6_mem_b2_b_59;
wire n_2456;
wire u3_mem_b3_b_152;
wire n_7769;
wire u6_mem_b2_b_58;
wire u10_mem_b1_b;
wire n_4403;
wire u6_mem_b2_b_34;
wire n_7774;
wire u6_mem_b2_b_54;
wire oc3_cfg_999;
wire n_8534;
wire n_1509;
wire n_7775;
wire u6_mem_b2_b_53;
wire n_8850;
wire n_4482;
wire n_7560;
wire n_8851;
wire n_4479;
wire n_7561;
wire n_3299;
wire n_8235;
wire u11_mem_b0_b_161;
wire n_10815;
wire n_9520;
wire n_9365;
wire n_6367;
wire n_6366;
wire n_9908;
wire n_9910;
wire n_9672;
wire n_4679;
wire n_9461;
wire n_8482;
wire n_9359;
wire n_9462;
wire n_8483;
wire n_8679;
wire n_9463;
wire n_8484;
wire n_9635;
wire n_9507;
wire n_9636;
wire n_9508;
wire n_9637;
wire n_9509;
wire n_9477;
wire n_4912;
wire n_3321;
wire n_3852;
wire u8_mem_b3_b_125;
wire n_1414;
wire n_4913;
wire u3_mem_b1_b_74;
wire n_2743;
wire n_4914;
wire u6_mem_b3_b_129;
wire n_3035;
wire n_4915;
wire u6_mem_b3_b_128;
wire n_4916;
wire u6_mem_b3_b_127;
wire n_4917;
wire u6_mem_b3_b_125;
wire n_3204;
wire n_4918;
wire u7_mem_b1_b_70;
wire n_2752;
wire n_3851;
wire u8_mem_b3_b_131;
wire n_6376;
wire n_6589;
wire u5_mem_b0_b_99;
wire n_9417;
wire n_6371;
wire n_6370;
wire n_10123;
wire n_6338;
wire n_6337;
wire n_10411;
wire n_6336;
wire n_10122;
wire n_6332;
wire n_6331;
wire n_9639;
wire u7_mem_b3_b;
wire n_8983;
wire n_9988;
wire n_313;
wire n_4399;
wire n_1990;
wire n_5065;
wire u4_mem_b3_b_129;
wire n_2992;
wire n_2486;
wire n_1067;
wire n_3864;
wire u8_mem_b3_b_124;
wire n_1478;
wire n_4397;
wire u8_mem_b1_b_82;
wire n_10367;
wire n_277;
wire n_4398;
wire n_2145;
wire i4_dout_600;
wire n_4811;
wire n_1507;
wire u3_mem_b3_b_126;
wire n_1517;
wire n_2379;
wire u3_mem_b3_b_149;
wire n_4396;
wire u8_mem_b2_b_49;
wire n_2164;
wire n_9872;
wire u10_din_tmp_43;
wire n_11119;
wire n_6515;
wire u11_mem_b1_b_130;
wire n_5533;
wire n_5813;
wire n_11447;
wire n_11448;
wire n_2338;
wire n_2455;
wire u8_mem_b2_b_34;
wire n_8473;
wire crac_din_694;
wire n_1047;
wire ic2_cfg;
wire n_8608;
wire n_6047;
wire n_3633;
wire oc5_int_set_718;
wire n_9573;
wire u11_mem_b3_b_73;
wire n_10834;
wire n_175;
wire n_8536;
wire n_3631;
wire n_3688;
wire n_8021;
wire u4_mem_b1_b_66;
wire n_12054;
wire n_1578;
wire n_6445;
wire n_1575;
wire n_6417;
wire n_1831;
wire n_1582;
wire n_1580;
wire n_1583;
wire n_190;
wire n_5508;
wire n_2521;
wire u10_din_tmp1;
wire u13_ints_r_b23_b;
wire n_9845;
wire n_12057;
wire n_2466;
wire n_3094;
wire n_6545;
wire n_8202;
wire n_8196;
wire n_4688;
wire n_8193;
wire n_4714;
wire n_8194;
wire n_8201;
wire wb_din_671;
wire oc5_cfg_1016;
wire n_8362;
wire n_8198;
wire n_8200;
wire n_8199;
wire n_930;
wire n_5535;
wire n_2445;
wire n_3398;
wire n_3404;
wire n_2244;
wire n_8192;
wire n_4711;
wire n_5498;
wire u11_mem_b3_b_84;
wire u11_din_tmp_52;
wire n_10112;
wire u11_wp_b2_b;
wire n_11852;
wire n_3921;
wire n_2475;
wire n_10267;
wire n_6496;
wire n_6495;
wire u3_mem_b0_b_96;
wire n_9366;
wire n_10289;
wire n_10250;
wire n_10290;
wire n_10287;
wire n_10288;
wire n_6648;
wire n_6647;
wire n_10295;
wire n_10308;
wire n_10296;
wire n_10291;
wire n_6538;
wire n_10293;
wire u7_mem_b1_b_90;
wire n_4121;
wire u7_mem_b2_b_59;
wire n_11729;
wire n_4123;
wire n_4124;
wire u7_mem_b1_b_88;
wire n_9629;
wire n_9579;
wire n_9472;
wire n_9471;
wire n_8644;
wire n_2181;
wire n_2059;
wire n_1472;
wire n_4117;
wire u7_mem_b1_b_84;
wire n_3920;
wire u10_din_tmp_51;
wire wb_din_684;
wire n_1363;
wire n_823;
wire n_434;
wire n_625;
wire n_10344;
wire n_9972;
wire n_1107;
wire n_1889;
wire n_908;
wire n_4703;
wire n_8581;
wire n_697;
wire n_6035;
wire n_1979;
wire u10_mem_b3_b_73;
wire n_8727;
wire n_1205;
wire n_1684;
wire u10_mem_b1_b_142;
wire n_1609;
wire u11_mem_b1_b_143;
wire n_9040;
wire n_1981;
wire u11_mem_b3_b_71;
wire n_10456;
wire n_1980;
wire n_1927;
wire u8_mem_b2_b_32;
wire n_909;
wire n_1982;
wire n_12583;
wire n_3922;
wire n_2335;
wire n_3683;
wire u6_mem_b0_b;
wire n_1983;
wire n_7207;
wire n_5906;
wire n_6156;
wire n_7120;
wire n_2352;
wire u8_mem_b2_b_46;
wire n_2366;
wire u15_crac_we_r;
wire n_2678;
wire n_7117;
wire n_5907;
wire n_5742;
wire u4_mem_b1_b_79;
wire n_8328;
wire n_11063;
wire n_7209;
wire n_6279;
wire n_5760;
wire n_7214;
wire n_7114;
wire n_5939;
wire n_5794;
wire n_7212;
wire n_8271;
wire n_4413;
wire n_8333;
wire n_7992;
wire n_7172;
wire n_5938;
wire n_5793;
wire n_3692;
wire u5_mem_b3_b_132;
wire n_9234;
wire n_4863;
wire n_7575;
wire n_7204;
wire n_6154;
wire n_3693;
wire u5_mem_b0_b_98;
wire n_7205;
wire n_6277;
wire n_3694;
wire wb_din_667;
wire n_3696;
wire u5_mem_b0_b_94;
wire n_6060;
wire n_6757;
wire n_116;
wire n_7011;
wire n_95;
wire n_6040;
wire n_4843;
wire n_796;
wire n_1255;
wire n_5964;
wire n_5637;
wire n_1443;
wire n_5636;
wire n_8355;
wire n_5121;
wire n_8357;
wire n_3690;
wire u5_mem_b0_b_95;
wire wb_din_665;
wire n_3790;
wire u4_mem_b0_b_95;
wire n_3765;
wire n_9516;
wire n_9361;
wire o9_empty;
wire o8_empty;
wire u10_mem_b0_b_176;
wire n_9515;
wire n_9360;
wire n_12502;
wire n_9460;
wire n_8183;
wire n_8678;
wire n_4571;
wire n_2385;
wire n_4954;
wire n_8057;
wire n_4231;
wire n_5282;
wire n_4230;
wire n_5287;
wire u13_ints_r_b21_b;
wire u8_mem_b2_b_54;
wire n_11446;
wire n_11445;
wire n_4310;
wire u4_mem_b2_b_40;
wire n_2016;
wire n_3436;
wire u3_mem_b0_b_115;
wire n_3986;
wire oc2_cfg_990;
wire n_7484;
wire u10_mem_b2_b_105;
wire n_10772;
wire n_4570;
wire n_3545;
wire n_2496;
wire n_4721;
wire u13_intm_r_b16_b;
wire u13_ints_r_b16_b;
wire n_8358;
wire n_5125;
wire n_8065;
wire n_1234;
wire n_512;
wire n_853;
wire n_3786;
wire n_515;
wire u26_ps_cnt_b4_b;
wire n_8794;
wire n_1558;
wire n_606;
wire u5_mem_b3_b_140;
wire u7_mem_b0_b_99;
wire n_9389;
wire n_3540;
wire u5_mem_b3_b_152;
wire n_3172;
wire n_9149;
wire n_9068;
wire n_3857;
wire n_8130;
wire n_4888;
wire u7_mem_b3_b_131;
wire n_3311;
wire n_835;
wire u3_mem_b1_b_81;
wire n_2670;
wire n_2705;
wire n_2846;
wire u8_mem_b1_b_68;
wire n_12301;
wire n_2672;
wire n_2770;
wire n_1969;
wire n_1965;
wire n_1966;
wire u3_mem_b2_b_54;
wire n_3330;
wire u5_mem_b2_b_29;
wire n_9261;
wire n_7073;
wire n_5682;
wire n_7077;
wire n_6191;
wire u3_mem_b0_b_112;
wire n_8842;
wire i3_dout_574;
wire n_4065;
wire n_11074;
wire u5_mem_b3_b_127;
wire n_9201;
wire n_3647;
wire u7_mem_b0_b_103;
wire n_8921;
wire n_2849;
wire n_11720;
wire u3_mem_b1_b_69;
wire n_12753;
wire n_7452;
wire u6_mem_b1_b_90;
wire n_9158;
wire n_9147;
wire u11_mem_b1_b_133;
wire u4_mem_b2_b_39;
wire n_8300;
wire n_10323;
wire n_3792;
wire n_8953;
wire n_10967;
wire u13_ints_r_b11_b;
wire n_11146;
wire n_9072;
wire n_4340;
wire n_8898;
wire n_7588;
wire u14_u6_en_out_l2;
wire n_1761;
wire n_6450;
wire n_4628;
wire n_2460;
wire n_1860;
wire n_6534;
wire n_1834;
wire n_6087;
wire n_1222;
wire n_2421;
wire n_3494;
wire n_1770;
wire n_6956;
wire n_1768;
wire n_6924;
wire n_1220;
wire n_1767;
wire n_1766;
wire n_1765;
wire n_6402;
wire n_6551;
wire n_1764;
wire n_6617;
wire n_1763;
wire n_6614;
wire n_9112;
wire n_4928;
wire n_9110;
wire n_7760;
wire n_9111;
wire n_7759;
wire ic2_cfg_1046;
wire n_8601;
wire n_9120;
wire n_9119;
wire n_4330;
wire n_7767;
wire n_9118;
wire n_4457;
wire n_7766;
wire n_9117;
wire n_4401;
wire n_9077;
wire n_7765;
wire n_9116;
wire n_7764;
wire n_7763;
wire n_9114;
wire n_4415;
wire n_7762;
wire n_9113;
wire n_4322;
wire n_7761;
wire n_3855;
wire u8_mem_b3_b_123;
wire n_2577;
wire n_4677;
wire n_2918;
wire n_2614;
wire u13_ints_r_b14_b;
wire n_935;
wire n_1019;
wire n_6056;
wire n_4805;
wire n_2938;
wire n_3406;
wire n_1406;
wire n_970;
wire n_6816;
wire n_837;
wire ic0_cfg_1026;
wire n_836;
wire oc3_cfg_995;
wire n_5633;
wire n_4101;
wire u9_mem_b3_b_62;
wire n_11174;
wire n_11021;
wire u5_mem_b2_b_36;
wire n_9239;
wire n_4058;
wire n_445;
wire n_868;
wire u8_mem_b2_b_40;
wire n_8885;
wire u11_mem_b2_b_93;
wire u9_mem_b0_b_170;
wire n_7446;
wire n_7378;
wire n_11888;
wire n_346;
wire n_345;
wire n_347;
wire n_343;
wire n_10029;
wire n_6089;
wire n_2499;
wire n_385;
wire n_12383;
wire n_551;
wire n_10028;
wire n_10027;
wire n_10024;
wire n_7448;
wire n_7379;
wire n_11887;
wire n_11711;
wire n_12204;
wire u6_mem_b0_b_95;
wire n_9079;
wire n_7496;
wire n_7870;
wire n_3154;
wire n_10335;
wire n_1798;
wire n_12640;
wire n_11666;
wire n_1796;
wire n_3158;
wire u8_mem_b1_b_88;
wire n_1795;
wire n_5749;
wire n_5181;
wire n_6093;
wire n_5747;
wire n_5748;
wire u13_intm_r_b13_b;
wire n_8516;
wire n_5753;
wire n_5195;
wire n_6094;
wire n_5452;
wire n_5453;
wire n_6118;
wire n_5744;
wire n_5745;
wire n_5182;
wire n_11563;
wire u9_mem_b2_b_104;
wire n_10279;
wire n_2441;
wire u3_mem_b3_b_142;
wire i6_dout_633;
wire n_4002;
wire u5_mem_b3_b_137;
wire n_9228;
wire n_4106;
wire n_5307;
wire n_8528;
wire n_8529;
wire n_3057;
wire n_11730;
wire n_3056;
wire n_2276;
wire u6_mem_b2_b_32;
wire n_4161;
wire n_1541;
wire u10_din_tmp_54;
wire n_9856;
wire n_3947;
wire u4_mem_b0_b_112;
wire n_9437;
wire n_6103;
wire n_4572;
wire n_5198;
wire u5_mem_b2_b_52;
wire n_9255;
wire u5_mem_b3_b_151;
wire n_4838;
wire n_3432;
wire n_4837;
wire n_5116;
wire n_7565;
wire n_7776;
wire n_8859;
wire n_4326;
wire n_7697;
wire n_8858;
wire n_4321;
wire n_7566;
wire n_8861;
wire n_4271;
wire n_7567;
wire n_8860;
wire n_4857;
wire n_7694;
wire n_8864;
wire n_7569;
wire crac_din_693;
wire n_1194;
wire n_3583;
wire u8_mem_b0_b_95;
wire n_4839;
wire n_10762;
wire n_3544;
wire u5_mem_b3_b_149;
wire n_8007;
wire u4_mem_b2_b_29;
wire n_8006;
wire u4_mem_b3_b_127;
wire n_7952;
wire u4_mem_b3_b_128;
wire u4_mem_b3_b_152;
wire u4_mem_b3_b_150;
wire n_8011;
wire u4_mem_b3_b_126;
wire n_7957;
wire u3_mem_b1_b_70;
wire n_8008;
wire u4_mem_b2_b_47;
wire n_12146;
wire n_12147;
wire i6_dout;
wire n_4032;
wire n_12142;
wire n_12143;
wire n_4086;
wire n_2599;
wire n_1814;
wire n_6790;
wire n_3731;
wire u5_mem_b0_b_106;
wire n_6803;
wire u5_mem_b2_b_51;
wire n_9256;
wire dma_req_o_b0_b;
wire n_11192;
wire n_10917;
wire u9_mem_b1_b_142;
wire n_10748;
wire n_6817;
wire n_6765;
wire n_3732;
wire n_10849;
wire u4_mem_b1_b_63;
wire n_8309;
wire n_3587;
wire n_9190;
wire n_3727;
wire n_9409;
wire n_3586;
wire u3_mem_b0_b_116;
wire n_3728;
wire u5_mem_b0_b_107;
wire n_3585;
wire u3_mem_b0_b_117;
wire wb_din_687;
wire n_7281;
wire n_6837;
wire n_2300;
wire n_840;
wire n_462;
wire n_6267;
wire n_7395;
wire n_7356;
wire n_8209;
wire n_5434;
wire n_10621;
wire u3_mem_b2_b_33;
wire n_8395;
wire n_10620;
wire n_10616;
wire n_10618;
wire n_10614;
wire n_6205;
wire n_6203;
wire n_10615;
wire n_4334;
wire n_2155;
wire n_4929;
wire n_2812;
wire n_4332;
wire n_7026;
wire n_7025;
wire n_1271;
wire u6_mem_b2_b_31;
wire n_1937;
wire n_4331;
wire u8_mem_b2_b_39;
wire n_2143;
wire u6_mem_b3_b;
wire n_4329;
wire u8_mem_b1_b_69;
wire n_2124;
wire n_4926;
wire n_3040;
wire n_7282;
wire n_6840;
wire n_2232;
wire u14_u1_en_out_l2;
wire n_9479;
wire n_12837;
wire n_6843;
wire n_9171;
wire n_7536;
wire n_3725;
wire u5_mem_b0_b_109;
wire n_7457;
wire n_6673;
wire n_615;
wire u11_mem_b2_b_107;
wire o6_status;
wire n_7296;
wire n_6737;
wire n_6693;
wire n_3719;
wire u5_mem_b0_b_111;
wire n_2126;
wire n_2129;
wire n_8748;
wire n_2764;
wire n_2689;
wire n_2132;
wire n_2131;
wire n_1920;
wire n_5325;
wire n_5298;
wire n_5326;
wire u11_mem_b1_b_144;
wire n_5309;
wire n_5334;
wire n_5333;
wire n_3948;
wire n_5336;
wire n_5335;
wire n_5405;
wire n_5337;
wire n_5338;
wire n_5296;
wire n_5327;
wire n_5321;
wire n_5329;
wire u11_mem_b1_b_141;
wire n_5313;
wire n_5331;
wire u10_mem_b2_b_117;
wire n_5330;
wire n_5332;
wire u11_mem_b1_b_140;
wire n_3722;
wire u5_mem_b0_b_110;
wire wb_din_680;
wire n_4428;
wire n_1992;
wire n_4948;
wire u6_mem_b1_b;
wire n_2675;
wire n_518;
wire ic2_cfg_1049;
wire n_4947;
wire n_2652;
wire u7_mem_b2_b_32;
wire n_2204;
wire n_3715;
wire u5_mem_b0_b_113;
wire n_4430;
wire u8_mem_b1_b_65;
wire n_2193;
wire n_6075;
wire u3_mem_b1_b_75;
wire n_8893;
wire n_4950;
wire n_3031;
wire n_11715;
wire n_11716;
wire n_1810;
wire n_2426;
wire n_1085;
wire u9_rp_b2_b;
wire n_737;
wire n_6977;
wire n_5529;
wire n_7063;
wire n_5896;
wire n_4949;
wire u7_mem_b3_b_136;
wire n_3501;
wire n_6951;
wire u9_mem_b3_b_73;
wire n_6882;
wire n_6881;
wire n_4614;
wire u9_din_tmp_48;
wire n_4616;
wire n_3932;
wire n_4350;
wire n_2292;
wire i3_dout_582;
wire n_4057;
wire n_1699;
wire n_1697;
wire n_5704;
wire n_3861;
wire u8_mem_b3_b_128;
wire n_4613;
wire n_12059;
wire n_2458;
wire n_3468;
wire n_1832;
wire n_4229;
wire n_3070;
wire n_1698;
wire n_6505;
wire n_2388;
wire n_3480;
wire n_1569;
wire n_3913;
wire u10_din_tmp_52;
wire n_12052;
wire n_4163;
wire n_3073;
wire n_8535;
wire oc0_cfg_965;
wire n_8537;
wire n_9056;
wire n_8543;
wire n_8545;
wire oc3_cfg_994;
wire n_8546;
wire n_1873;
wire n_8548;
wire n_8549;
wire n_3987;
wire n_8551;
wire n_10262;
wire n_6621;
wire n_6620;
wire n_10263;
wire n_6926;
wire n_10277;
wire n_10264;
wire n_6629;
wire n_6628;
wire n_10266;
wire n_6929;
wire n_6928;
wire n_10651;
wire n_6624;
wire n_6623;
wire n_10268;
wire n_6901;
wire n_11032;
wire n_8781;
wire n_10259;
wire n_6615;
wire n_10261;
wire n_6619;
wire n_6922;
wire u9_mem_b3_b_72;
wire n_4113;
wire n_11856;
wire n_12721;
wire n_2915;
wire u8_mem_b1_b_86;
wire n_2913;
wire u3_mem_b2_b_49;
wire n_1211;
wire u11_mem_b2_b_100;
wire n_1214;
wire u11_mem_b2_b_110;
wire n_10870;
wire n_438;
wire n_12332;
wire u11_mem_b1_b_131;
wire n_10843;
wire n_3606;
wire n_8980;
wire n_7650;
wire n_2376;
wire u6_mem_b3_b_124;
wire n_12622;
wire u9_mem_b2_b_105;
wire u26_cnt_b1_b;
wire n_9493;
wire n_8985;
wire n_4294;
wire n_7655;
wire n_9703;
wire n_9421;
wire n_8556;
wire n_3608;
wire n_12802;
wire n_485;
wire n_422;
wire n_3526;
wire u5_mem_b3_b_141;
wire n_11135;
wire u6_mem_b0_b_99;
wire n_9402;
wire u9_mem_b0_b_162;
wire n_10170;
wire o8_status_1002;
wire i6_dout_637;
wire o7_status_992;
wire i6_dout_638;
wire i3_dout_576;
wire o6_status_982;
wire n_6683;
wire i3_dout_571;
wire n_7161;
wire o4_status_972;
wire n_6680;
wire i6_dout_626;
wire i3_dout_564;
wire n_2115;
wire n_2790;
wire i6_dout_635;
wire i3_dout_573;
wire n_7113;
wire n_5892;
wire u13_ints_r_b1_b;
wire o9_status_1012;
wire n_749;
wire ic2_int_set_724;
wire n_221;
wire n_699;
wire n_1083;
wire n_523;
wire ic1_cfg_1039;
wire n_10820;
wire n_9903;
wire u3_mem_b3_b_140;
wire n_8376;
wire n_11529;
wire n_9413;
wire n_3313;
wire n_125;
wire n_5524;
wire n_2700;
wire u4_mem_b0_b_114;
wire n_11472;
wire n_12261;
wire u7_mem_b3_b_146;
wire n_3426;
wire n_2676;
wire n_2736;
wire n_2644;
wire n_3428;
wire n_4834;
wire n_1377;
wire u6_rp_b3_b;
wire n_11040;
wire n_8594;
wire u2_to_cnt_b0_b;
wire n_8413;
wire n_1588;
wire n_6498;
wire n_11152;
wire n_6053;
wire n_12639;
wire n_11494;
wire u5_mem_b2_b;
wire n_1600;
wire n_1599;
wire n_8756;
wire n_3664;
wire n_7505;
wire n_9405;
wire u6_mem_b0_b_94;
wire n_3648;
wire n_3663;
wire n_8755;
wire u6_mem_b0_b_96;
wire n_3652;
wire n_8759;
wire u6_mem_b0_b_120;
wire n_3667;
wire n_8758;
wire n_3628;
wire n_9406;
wire u6_mem_b0_b_121;
wire n_3666;
wire n_3658;
wire n_3660;
wire n_1596;
wire n_1595;
wire u4_mem_b2_b_56;
wire n_8278;
wire u3_mem_b3_b_131;
wire n_8388;
wire n_188;
wire n_1662;
wire n_6363;
wire u9_mem_b2_b_93;
wire n_7528;
wire n_568;
wire n_936;
wire u8_mem_b0_b_118;
wire n_9378;
wire n_1592;
wire n_1591;
wire crac_din_702;
wire n_1029;
wire n_4666;
wire n_5292;
wire n_6594;
wire n_2400;
wire u8_mem_b3_b_150;
wire n_4964;
wire n_2793;
wire n_4963;
wire n_4615;
wire u9_din_tmp_47;
wire n_4349;
wire n_4965;
wire u5_mem_b3_b_130;
wire n_4611;
wire n_2374;
wire n_2863;
wire n_4967;
wire u6_mem_b1_b_77;
wire n_5019;
wire n_2809;
wire n_4966;
wire u5_mem_b3_b_129;
wire n_5224;
wire n_4109;
wire n_3134;
wire n_1696;
wire n_6909;
wire n_3860;
wire u8_mem_b3_b_151;
wire n_4962;
wire u7_mem_b3_b_137;
wire n_3455;
wire n_9195;
wire n_4346;
wire n_7835;
wire n_9193;
wire n_3850;
wire n_7727;
wire n_9197;
wire n_3858;
wire n_7837;
wire n_9196;
wire n_7596;
wire n_7830;
wire n_9189;
wire n_4933;
wire n_7828;
wire n_9192;
wire n_7832;
wire n_9191;
wire n_4930;
wire n_7831;
wire n_9188;
wire n_4946;
wire n_7827;
wire n_4938;
wire n_7825;
wire n_8870;
wire n_4872;
wire n_7572;
wire u7_mem_b3_b_139;
wire n_5516;
wire u10_mem_b3_b_79;
wire n_3959;
wire n_4745;
wire u8_mem_b2_b_37;
wire n_8469;
wire n_3960;
wire u10_mem_b1_b_141;
wire n_10671;
wire n_4278;
wire n_7573;
wire n_3961;
wire n_4085;
wire n_4747;
wire n_4667;
wire n_3137;
wire n_4669;
wire n_3138;
wire n_4668;
wire n_3275;
wire u7_mem_b3_b_130;
wire n_8872;
wire n_4270;
wire n_7580;
wire n_1525;
wire n_1055;
wire n_1104;
wire n_680;
wire u9_mem_b2_b_113;
wire n_8189;
wire n_9855;
wire n_6408;
wire u10_mem_b1_b_124;
wire n_1620;
wire u11_mem_b0_b_172;
wire n_2526;
wire n_5945;
wire u3_wp_b0_b;
wire n_418;
wire oc4_cfg;
wire u11_mem_b2_b_98;
wire n_508;
wire n_8286;
wire n_1167;
wire n_12627;
wire n_4175;
wire n_4191;
wire n_2993;
wire n_1339;
wire n_12807;
wire u5_mem_b1_b_65;
wire n_10006;
wire n_5514;
wire n_10005;
wire u10_mem_b3_b_69;
wire n_10229;
wire u5_wp_b1_b;
wire n_10011;
wire n_5520;
wire n_10009;
wire n_5363;
wire n_10008;
wire n_5518;
wire n_10007;
wire n_9759;
wire n_9608;
wire n_9454;
wire n_10013;
wire n_5577;
wire n_10012;
wire n_669;
wire n_11737;
wire n_7402;
wire n_10769;
wire n_4793;
wire n_10450;
wire n_10079;
wire n_10770;
wire n_5380;
wire n_10080;
wire n_1106;
wire o9_status;
wire n_847;
wire o8_status;
wire n_10771;
wire n_5425;
wire n_10082;
wire n_5426;
wire n_10679;
wire n_10084;
wire n_9644;
wire o4_status;
wire n_9606;
wire n_7408;
wire o6_we;
wire n_9286;
wire n_9583;
wire n_1391;
wire n_5421;
wire n_4036;
wire n_5576;
wire n_4819;
wire n_5578;
wire n_4820;
wire n_4075;
wire n_4074;
wire n_1813;
wire n_6088;
wire n_5569;
wire n_6090;
wire n_5570;
wire n_5734;
wire u9_mem_b2_b_106;
wire n_5733;
wire n_5735;
wire n_5736;
wire n_5423;
wire u10_mem_b1_b_137;
wire n_5422;
wire n_5737;
wire u9_mem_b1_b_136;
wire n_4690;
wire n_11894;
wire n_9717;
wire n_9666;
wire u9_mem_b2_b_114;
wire n_6528;
wire u9_mem_b1_b_133;
wire n_6625;
wire u11_mem_b3_b_63;
wire u10_mem_b2_b_118;
wire n_10733;
wire u9_mem_b0_b;
wire n_10176;
wire n_8879;
wire n_4495;
wire n_7577;
wire n_8311;
wire n_8086;
wire u3_mem_b3_b_146;
wire n_1379;
wire n_4873;
wire n_8387;
wire n_8102;
wire n_8084;
wire u3_mem_b3_b_148;
wire n_3565;
wire n_8083;
wire n_8081;
wire u3_mem_b3_b_150;
wire i4_dout_609;
wire n_5393;
wire n_8082;
wire n_10321;
wire n_6665;
wire n_6664;
wire n_10319;
wire n_6663;
wire n_6662;
wire n_10318;
wire n_6661;
wire n_6660;
wire n_10317;
wire n_6034;
wire n_10316;
wire n_6031;
wire n_5137;
wire n_8095;
wire n_10314;
wire n_6957;
wire n_10313;
wire n_6657;
wire n_6656;
wire n_10311;
wire n_6552;
wire n_10310;
wire n_6541;
wire n_8080;
wire n_8079;
wire n_8078;
wire n_1362;
wire u7_mem_b3_b_122;
wire n_5506;
wire n_9411;
wire n_7756;
wire u6_mem_b3_b_133;
wire n_8880;
wire n_4864;
wire n_7578;
wire n_4866;
wire n_7585;
wire n_8892;
wire n_4328;
wire n_7584;
wire n_8890;
wire n_4273;
wire n_7583;
wire n_4865;
wire n_7791;
wire u6_mem_b2_b_37;
wire n_8883;
wire n_8125;
wire n_3530;
wire u4_mem_b3_b_144;
wire n_3556;
wire n_7673;
wire n_2273;
wire n_4155;
wire n_2272;
wire u6_mem_b2_b_33;
wire n_3045;
wire u3_mem_b1_b_88;
wire n_12819;
wire u6_mem_b2_b_29;
wire n_3236;
wire n_12822;
wire u6_mem_b1_b_62;
wire n_12821;
wire n_3044;
wire n_3043;
wire n_8361;
wire n_5130;
wire n_7619;
wire n_8360;
wire n_4953;
wire n_7974;
wire u4_mem_b3_b_138;
wire n_7973;
wire u4_mem_b3_b_139;
wire n_7972;
wire n_7971;
wire u4_mem_b3_b_122;
wire n_681;
wire n_8354;
wire n_5124;
wire n_8074;
wire n_8353;
wire n_4908;
wire n_8073;
wire n_7515;
wire n_12124;
wire n_12120;
wire n_12121;
wire u3_rp_b1_b;
wire n_11162;
wire u11_mem_b1_b_122;
wire n_10551;
wire n_9084;
wire o3_we;
wire n_7028;
wire u10_mem_b0_b_161;
wire n_10451;
wire n_10710;
wire n_7437;
wire crac_out_863;
wire n_8634;
wire u6_mem_b3_b_142;
wire n_3167;
wire u9_din_tmp_50;
wire n_9770;
wire u10_mem_b2_b_92;
wire n_5988;
wire u11_mem_b1_b_135;
wire n_795;
wire n_8715;
wire n_141;
wire n_11748;
wire n_12453;
wire n_10599;
wire n_10601;
wire n_10592;
wire n_11634;
wire n_11096;
wire n_8182;
wire n_10595;
wire n_11616;
wire n_11614;
wire n_11891;
wire n_9668;
wire n_11889;
wire n_12501;
wire n_3755;
wire u4_mem_b0_b_96;
wire n_4935;
wire n_2811;
wire n_4936;
wire n_2750;
wire u8_mem_b2_b_56;
wire n_1989;
wire n_4435;
wire n_2188;
wire n_4440;
wire u9_din_tmp_42;
wire n_9779;
wire n_4942;
wire u6_mem_b1_b_79;
wire n_2664;
wire n_4943;
wire u6_mem_b1_b_60;
wire n_2709;
wire n_4937;
wire n_2824;
wire n_2680;
wire n_4939;
wire u6_mem_b1_b_87;
wire n_2826;
wire u11_mem_b1_b_129;
wire n_10561;
wire n_11893;
wire n_11777;
wire u11_mem_b0_b_155;
wire n_10420;
wire n_2527;
wire n_11919;
wire n_11908;
wire n_11914;
wire n_2107;
wire n_11504;
wire n_2113;
wire n_2111;
wire n_2110;
wire n_2757;
wire n_2109;
wire n_2114;
wire n_2108;
wire n_2071;
wire n_8588;
wire n_4713;
wire u11_rp_b1_b;
wire n_7375;
wire n_10535;
wire n_3759;
wire u4_mem_b0_b_121;
wire n_12520;
wire n_12516;
wire n_12517;
wire n_12604;
wire n_1320;
wire n_1084;
wire n_532;
wire n_12330;
wire n_10306;
wire i3_dout_569;
wire n_4041;
wire n_1121;
wire n_3517;
wire n_12839;
wire n_4249;
wire u6_mem_b1_b_76;
wire n_1432;
wire n_12752;
wire n_11719;
wire u3_mem_b0_b_100;
wire n_8261;
wire n_3519;
wire n_818;
wire u26_ps_cnt_b0_b;
wire n_3520;
wire n_1629;
wire n_1317;
wire n_6565;
wire n_7927;
wire n_976;
wire n_498;
wire n_1638;
wire n_6500;
wire n_1639;
wire n_6654;
wire n_5212;
wire n_4183;
wire n_1637;
wire n_6454;
wire n_6413;
wire n_1635;
wire n_1634;
wire n_3588;
wire n_1631;
wire n_4581;
wire n_2258;
wire n_8570;
wire oc1_cfg_975;
wire n_3524;
wire u3_mem_b0_b_111;
wire n_3171;
wire u7_mem_b0_b_98;
wire n_8584;
wire n_4708;
wire n_8586;
wire n_4710;
wire n_4699;
wire n_8575;
wire n_8577;
wire ic0_cfg_1030;
wire n_8571;
wire n_8573;
wire ic1_cfg_1034;
wire n_10243;
wire n_6897;
wire n_6895;
wire n_10244;
wire n_6022;
wire n_10241;
wire n_6887;
wire n_10242;
wire n_6914;
wire n_10600;
wire n_6019;
wire n_6018;
wire n_10239;
wire n_6910;
wire n_10236;
wire n_6907;
wire n_10233;
wire n_6603;
wire n_6601;
wire n_10234;
wire n_6006;
wire n_9584;
wire o3_status;
wire n_9556;
wire n_2433;
wire u8_mem_b3_b_140;
wire n_3596;
wire in_valid_s1;
wire n_9643;
wire u6_mem_b1_b_67;
wire n_4518;
wire n_4520;
wire u3_mem_b2_b_57;
wire n_2263;
wire n_6085;
wire n_7187;
wire n_6785;
wire n_7184;
wire n_6069;
wire n_5842;
wire n_1907;
wire n_5551;
wire n_5848;
wire o9_we;
wire n_7023;
wire n_5549;
wire n_5846;
wire n_5854;
wire n_6787;
wire n_5552;
wire n_5852;
wire n_6074;
wire n_5850;
wire n_4522;
wire n_1971;
wire n_2225;
wire n_3595;
wire u3_mem_b0_b_110;
wire n_12838;
wire n_4797;
wire n_4385;
wire n_6096;
wire n_5210;
wire n_4592;
wire n_9307;
wire n_9288;
wire n_9202;
wire n_9230;
wire n_9205;
wire n_4794;
wire u9_mem_b1_b_140;
wire n_3993;
wire n_3992;
wire n_4591;
wire n_3274;
wire n_2982;
wire n_2540;
wire n_2539;
wire n_2538;
wire n_1527;
wire n_1528;
wire u7_mem_b3_b_128;
wire n_5628;
wire u2_sync_resume;
wire n_7371;
wire n_7141;
wire n_6674;
wire n_7331;
wire n_7487;
wire n_7330;
wire n_7486;
wire n_6699;
wire n_7336;
wire n_7143;
wire n_7112;
wire n_7335;
wire n_6685;
wire n_7333;
wire n_7483;
wire n_6690;
wire n_7332;
wire n_7482;
wire n_6697;
wire n_9645;
wire n_571;
wire n_941;
wire u6_wp_b1_b;
wire n_9766;
wire n_1176;
wire n_2917;
wire u3_mem_b0_b_92;
wire n_10204;
wire n_7247;
wire n_7087;
wire n_8640;
wire u13_intm_r_b3_b;
wire n_8493;
wire n_8456;
wire i6_dout_644;
wire n_4021;
wire n_11044;
wire u7_mem_b2_b_44;
wire n_4753;
wire n_1870;
wire oc2_int_set;
wire n_9849;
wire n_1875;
wire n_2922;
wire n_12844;
wire u8_mem_b0_b_92;
wire n_1493;
wire u8_mem_b0_b_106;
wire n_691;
wire n_4223;
wire u7_mem_b1_b_87;
wire n_1453;
wire n_2435;
wire n_8975;
wire n_728;
wire u13_intm_r_b5_b;
wire u13_ints_r_b5_b;
wire u13_intm_r_b6_b;
wire u13_ints_r_b6_b;
wire n_8770;
wire u6_mem_b0_b_110;
wire n_3609;
wire n_8772;
wire u6_mem_b0_b_91;
wire n_3630;
wire n_8773;
wire n_8775;
wire n_9412;
wire n_8776;
wire n_9414;
wire n_8778;
wire u3_mem_b2_b_42;
wire n_9318;
wire u10_mem_b0_b_151;
wire n_10412;
wire u10_mem_b0_b_158;
wire n_12135;
wire n_12131;
wire n_12132;
wire n_11182;
wire n_11158;
wire u16_u3_dma_req_r1;
wire n_11172;
wire n_11124;
wire u16_u2_dma_req_r1;
wire n_11183;
wire n_11159;
wire u16_u1_dma_req_r1;
wire n_11173;
wire n_11125;
wire u16_u0_dma_req_r1;
wire n_4987;
wire n_2975;
wire n_4986;
wire n_5000;
wire n_3449;
wire n_4985;
wire u5_mem_b3_b_142;
wire n_3053;
wire n_4984;
wire n_3131;
wire n_4983;
wire u5_mem_b3_b_144;
wire n_3129;
wire n_9300;
wire n_4981;
wire u5_mem_b3_b_146;
wire n_3001;
wire n_4980;
wire n_3006;
wire n_6783;
wire n_11515;
wire n_2414;
wire n_4804;
wire n_5413;
wire n_4803;
wire n_5410;
wire n_6184;
wire n_3135;
wire n_3405;
wire n_1378;
wire n_3808;
wire u3_mem_b0_b;
wire n_5893;
wire n_3355;
wire n_2861;
wire n_2295;
wire n_2381;
wire n_5668;
wire n_7801;
wire n_9157;
wire n_7800;
wire n_1534;
wire u5_mem_b3_b_134;
wire n_9166;
wire n_7806;
wire n_9164;
wire n_7804;
wire n_9162;
wire n_7803;
wire n_7802;
wire n_4940;
wire n_7810;
wire n_9169;
wire n_5008;
wire n_7809;
wire n_9168;
wire n_5011;
wire n_7808;
wire n_9167;
wire n_5020;
wire n_7807;
wire oc0_int_set_707;
wire n_10907;
wire n_9596;
wire n_1535;
wire u9_mem_b1_b_121;
wire n_10299;
wire u12_re2;
wire u4_mem_b0_b_98;
wire n_8811;
wire n_4701;
wire n_454;
wire u11_mem_b0_b_178;
wire n_9175;
wire u5_mem_b1_b_88;
wire n_9289;
wire n_6220;
wire n_6221;
wire n_6153;
wire n_5438;
wire n_2566;
wire n_5830;
wire n_5829;
wire n_1772;
wire n_5834;
wire n_6782;
wire n_6781;
wire n_6780;
wire n_10652;
wire n_6029;
wire n_6028;
wire u10_mem_b1_b_131;
wire n_10211;
wire n_601;
wire u3_rp_b2_b;
wire n_6581;
wire u9_mem_b3_b_71;
wire u10_mem_b0_b_150;
wire u9_mem_b3_b_82;
wire u9_mem_b1_b_139;
wire n_63;
wire u9_mem_b2_b_117;
wire u11_mem_b0_b_177;
wire n_10433;
wire n_984;
wire n_1356;
wire n_9614;
wire n_1101;
wire n_5630;
wire n_5629;
wire n_2611;
wire n_1188;
wire n_1160;
wire u10_mem_b0_b_175;
wire n_5408;
wire u10_mem_b1_b_136;
wire n_5418;
wire n_1821;
wire u26_cnt_b2_b;
wire n_5406;
wire n_1820;
wire n_2612;
wire n_786;
wire n_1164;
wire n_4072;
wire n_1438;
wire n_5703;
wire n_6224;
wire u10_mem_b2_b_88;
wire u11_mem_b0_b_169;
wire n_10445;
wire i4_dout_613;
wire n_5390;
wire n_8931;
wire n_10892;
wire u4_mem_b3_b_141;
wire n_9343;
wire n_4754;
wire n_9995;
wire n_10750;
wire n_10059;
wire n_10751;
wire n_10060;
wire n_5342;
wire n_10058;
wire n_10753;
wire n_4790;
wire n_10062;
wire n_10754;
wire n_4791;
wire n_10063;
wire n_10755;
wire n_5731;
wire n_9991;
wire n_11722;
wire n_3183;
wire n_10055;
wire n_10744;
wire n_4750;
wire n_10056;
wire n_8918;
wire n_7601;
wire u6_mem_b1_b_71;
wire n_7822;
wire n_7821;
wire n_7824;
wire u6_mem_b1_b_74;
wire n_7823;
wire u6_mem_b1_b_75;
wire n_7819;
wire n_7818;
wire n_8867;
wire n_6438;
wire n_6437;
wire n_10508;
wire n_10501;
wire n_6446;
wire n_10190;
wire n_10187;
wire n_10197;
wire n_6452;
wire n_502;
wire n_10194;
wire n_5975;
wire n_5974;
wire n_10489;
wire n_10838;
wire n_6531;
wire n_6530;
wire n_732;
wire u10_mem_b2_b_104;
wire n_713;
wire u26_cnt_b0_b;
wire n_2314;
wire u4_mem_b2_b_30;
wire n_3223;
wire n_12842;
wire n_12041;
wire u5_mem_b2_b_43;
wire n_12364;
wire n_4494;
wire n_7579;
wire n_4460;
wire n_8039;
wire n_7755;
wire u6_mem_b3_b_134;
wire u4_mem_b2_b_31;
wire n_8272;
wire u9_mem_b3_b_65;
wire n_8169;
wire i6_dout_641;
wire i4_dout_610;
wire n_1851;
wire n_8171;
wire u8_mem_b2_b_35;
wire u10_mem_b2_b_96;
wire u6_mem_b1_b_63;
wire n_9156;
wire n_8334;
wire n_4464;
wire n_8336;
wire n_4475;
wire n_2589;
wire n_8439;
wire n_1429;
wire n_12624;
wire n_12630;
wire n_12632;
wire u6_mem_b2_b_36;
wire n_10406;
wire n_10087;
wire n_8886;
wire n_7805;
wire n_4344;
wire n_7582;
wire n_7757;
wire n_9466;
wire oc5_cfg_1019;
wire n_4420;
wire n_4421;
wire u4_mem_b2_b_55;
wire n_1970;
wire n_5110;
wire n_4422;
wire u4_mem_b2_b_54;
wire n_2048;
wire n_4423;
wire u4_mem_b2_b_53;
wire n_2484;
wire u7_mem_b2_b_40;
wire n_1994;
wire n_4425;
wire n_1998;
wire n_4426;
wire n_2100;
wire n_3348;
wire n_4419;
wire u4_mem_b2_b_57;
wire n_2024;
wire n_5109;
wire n_3507;
wire n_6268;
wire n_7048;
wire n_5902;
wire n_2226;
wire n_5904;
wire n_5859;
wire n_3559;
wire n_2095;
wire n_2094;
wire n_2093;
wire n_2091;
wire n_5903;
wire u6_mem_b1_b_84;
wire u5_mem_b3_b_150;
wire n_9210;
wire n_2746;
wire n_1082;
wire n_5021;
wire n_5022;
wire n_2806;
wire n_5018;
wire u5_mem_b1_b_89;
wire n_2828;
wire u6_mem_b1_b_86;
wire n_5016;
wire n_2800;
wire n_5017;
wire u5_mem_b1_b_90;
wire n_2719;
wire n_5014;
wire u5_mem_b1_b_64;
wire n_5015;
wire u5_mem_b1_b_63;
wire n_2967;
wire n_5012;
wire u5_mem_b1_b_66;
wire n_2835;
wire n_10377;
wire n_11797;
wire ic0_int_set_720;
wire n_5173;
wire n_2935;
wire resume_req;
wire n_7970;
wire oc5_int_set_717;
wire n_5631;
wire n_4100;
wire n_5170;
wire n_2870;
wire n_9275;
wire n_5010;
wire n_7907;
wire n_8363;
wire n_5066;
wire n_4698;
wire oc4_cfg_1010;
wire n_5260;
wire u13_intm_r_b7_b;
wire crac_din_698;
wire n_4697;
wire n_4704;
wire n_5263;
wire crac_din_696;
wire n_8784;
wire n_5261;
wire crac_din_697;
wire n_6000;
wire n_1602;
wire n_122;
wire n_5522;
wire n_4695;
wire oc5_cfg_1014;
wire n_5256;
wire u13_intm_r_b9_b;
wire crac_din_700;
wire n_8624;
wire n_8626;
wire crac_out_876;
wire n_8627;
wire crac_out_867;
wire n_8628;
wire crac_out_866;
wire n_8616;
wire n_4734;
wire n_8618;
wire n_4736;
wire n_8622;
wire n_4738;
wire n_8610;
wire ic1_cfg_1040;
wire u7_mem_b2_b_36;
wire n_1560;
wire n_5944;
wire n_657;
wire n_5942;
wire n_5901;
wire n_4841;
wire n_799;
wire n_1788;
wire n_4091;
wire n_1418;
wire n_1267;
wire n_4090;
wire n_1422;
wire n_1265;
wire n_6330;
wire n_6328;
wire n_10844;
wire n_6516;
wire n_6518;
wire n_6517;
wire u11_mem_b1_b_146;
wire n_10884;
wire n_3534;
wire n_3546;
wire n_10217;
wire n_6564;
wire n_6562;
wire n_10219;
wire n_6567;
wire n_10220;
wire n_6571;
wire n_6569;
wire n_10221;
wire n_6574;
wire n_6572;
wire n_10562;
wire n_6520;
wire n_6519;
wire n_10563;
wire n_6523;
wire n_10564;
wire n_6001;
wire n_10216;
wire n_6004;
wire n_6002;
wire n_8649;
wire u7_mem_b2_b;
wire u11_mem_b0_b_164;
wire n_10813;
wire n_1420;
wire n_11851;
wire n_3417;
wire n_11585;
wire n_2191;
wire u10_mem_b2_b_102;
wire n_1225;
wire n_621;
wire n_9427;
wire n_1028;
wire n_8318;
wire n_7414;
wire n_11892;
wire n_2742;
wire n_2685;
wire n_2154;
wire n_7111;
wire n_5268;
wire n_4749;
wire n_5361;
wire u10_mem_b1_b_135;
wire n_2683;
wire n_5613;
wire n_4830;
wire n_2622;
wire n_6755;
wire n_5612;
wire n_4835;
wire n_1918;
wire n_4082;
wire n_8565;
wire n_942;
wire n_785;
wire u5_rp_b3_b;
wire n_5444;
wire n_4084;
wire n_731;
wire n_577;
wire u10_mem_b3_b_60;
wire n_3334;
wire n_1434;
wire i4_dout_597;
wire n_4813;
wire n_2403;
wire n_1178;
wire n_714;
wire n_12274;
wire u3_mem_b2_b_50;
wire n_8406;
wire n_11033;
wire u8_mem_b1_b_81;
wire n_2350;
wire n_1460;
wire n_3400;
wire n_3401;
wire u4_mem_b2_b_58;
wire n_12831;
wire u3_mem_b1_b;
wire u4_mem_b1_b_80;
wire n_12265;
wire u10_mem_b3_b_61;
wire n_6852;
wire u9_mem_b0_b_154;
wire n_2950;
wire n_4218;
wire u10_mem_b3_b_78;
wire n_6607;
wire u10_mem_b2_b_94;
wire n_1881;
wire u8_mem_b3_b_127;
wire n_9846;
wire u11_mem_b3_b_87;
wire n_4257;
wire n_4258;
wire n_5347;
wire u9_mem_b3_b_84;
wire n_11025;
wire n_9422;
wire u5_mem_b0_b_114;
wire n_3714;
wire u11_din_tmp_53;
wire n_10111;
wire n_8789;
wire n_8791;
wire n_8787;
wire n_268;
wire dma_req_o_b4_b;
wire u11_mem_b0_b_151;
wire n_11036;
wire u8_mem_b1_b_85;
wire n_8916;
wire n_11070;
wire n_8694;
wire n_8160;
wire u13_intm_r_b23_b;
wire n_8505;
wire n_1724;
wire n_11191;
wire n_105;
wire n_11194;
wire n_278;
wire n_271;
wire n_11189;
wire n_284;
wire n_11170;
wire n_11190;
wire n_11171;
wire n_9302;
wire n_3552;
wire n_5530;
wire n_5807;
wire n_11455;
wire n_11456;
wire n_1867;
wire n_2390;
wire n_5001;
wire u5_mem_b3_b_131;
wire n_4999;
wire n_2929;
wire n_6070;
wire n_4226;
wire n_2333;
wire n_1376;
wire n_5531;
wire n_5815;
wire n_11457;
wire n_11458;
wire n_2128;
wire n_1892;
wire n_5673;
wire n_11895;
wire n_5002;
wire u5_mem_b3_b;
wire n_3023;
wire n_7456;
wire u5_mem_b3_b_145;
wire n_9217;
wire i4_dout_616;
wire n_5386;
wire n_9675;
wire n_9308;
wire dma_req_o_b1_b;
wire n_1727;
wire u11_mem_b1_b_120;
wire u3_mem_b1_b_86;
wire n_8347;
wire oc4_int_set_715;
wire n_96;
wire u10_mem_b1_b_143;
wire n_11030;
wire n_2142;
wire n_2147;
wire n_2149;
wire n_2151;
wire u10_mem_b1_b_126;
wire n_10179;
wire n_2153;
wire n_5596;
wire n_829;
wire n_11149;
wire n_1804;
wire n_5597;
wire n_844;
wire i3_status;
wire n_6232;
wire n_5847;
wire n_734;
wire n_5439;
wire n_807;
wire i6_status;
wire n_8338;
wire u9_mem_b3_b_61;
wire n_2956;
wire u9_mem_b2_b_88;
wire n_12366;
wire n_6419;
wire n_12376;
wire n_12375;
wire u9_mem_b2_b_94;
wire n_2488;
wire n_411;
wire ic0_cfg;
wire n_12614;
wire u9_mem_b0_b_173;
wire n_10159;
wire u5_mem_b2_b_41;
wire n_9269;
wire u5_mem_b1_b_70;
wire n_9315;
wire n_5398;
wire n_4070;
wire n_5396;
wire n_449;
wire n_4088;
wire n_2500;
wire u9_mem_b0_b_178;
wire u11_mem_b1_b_126;
wire n_6890;
wire u9_mem_b3_b_59;
wire n_11017;
wire n_1059;
wire n_8947;
wire n_3777;
wire n_12165;
wire u6_mem_b2_b_38;
wire u10_mem_b2_b_99;
wire n_10322;
wire out_slt9;
wire n_11102;
wire i6_full;
wire n_9030;
wire n_11631;
wire n_11632;
wire n_11018;
wire n_11639;
wire n_11640;
wire n_9474;
wire n_7295;
wire n_7526;
wire n_8915;
wire n_11016;
wire n_11641;
wire n_11642;
wire n_9526;
wire n_7387;
wire n_9446;
wire n_9885;
wire n_10787;
wire n_9836;
wire n_9691;
wire n_10338;
wire n_10900;
wire n_10337;
wire n_9961;
wire n_11439;
wire u5_mem_b2_b_31;
wire n_3192;
wire n_1483;
wire n_11444;
wire n_3199;
wire n_9626;
wire n_12148;
wire n_1604;
wire n_7797;
wire n_8936;
wire n_4287;
wire n_8941;
wire n_4412;
wire n_7982;
wire n_8940;
wire n_7615;
wire n_8939;
wire n_4288;
wire n_4885;
wire n_8951;
wire n_7623;
wire n_8946;
wire n_4956;
wire n_7622;
wire n_8945;
wire n_7621;
wire n_8425;
wire n_6027;
wire n_6026;
wire n_10185;
wire n_6527;
wire n_6526;
wire n_6414;
wire n_10184;
wire n_6416;
wire n_6415;
wire n_10183;
wire n_6543;
wire n_6542;
wire n_10182;
wire n_6412;
wire n_6411;
wire n_10454;
wire n_6525;
wire n_6524;
wire n_10181;
wire n_6409;
wire n_10453;
wire n_6418;
wire n_8274;
wire n_757;
wire u8_rp_b1_b;
wire n_11466;
wire u8_mem_b2_b_47;
wire n_6042;
wire n_1300;
wire n_7945;
wire n_9780;
wire n_8234;
wire u11_mem_b0_b_154;
wire n_7514;
wire n_7595;
wire u8_mem_b1_b_61;
wire n_6702;
wire i6_dout_640;
wire i3_dout_578;
wire i6_dout_647;
wire i6_dout_646;
wire i3_dout_584;
wire n_6706;
wire i3_dout;
wire n_5450;
wire n_6703;
wire i6_dout_639;
wire i3_dout_577;
wire i6_dout_651;
wire i3_dout_589;
wire i6_dout_648;
wire i3_dout_586;
wire n_10939;
wire u11_mem_b3_b_59;
wire u5_mem_b2_b_35;
wire n_9240;
wire n_4059;
wire n_1297;
wire n_834;
wire n_744;
wire u4_wp_b0_b;
wire n_12609;
wire n_12608;
wire n_12606;
wire n_5571;
wire n_6995;
wire n_5862;
wire n_12602;
wire n_12601;
wire n_5867;
wire n_12603;
wire n_242;
wire n_12605;
wire n_2135;
wire n_6845;
wire u9_mem_b0_b_158;
wire n_632;
wire n_8513;
wire n_5886;
wire n_12030;
wire n_3260;
wire n_12031;
wire n_1340;
wire n_1274;
wire n_576;
wire n_442;
wire n_726;
wire n_8319;
wire n_5720;
wire n_5566;
wire n_3270;
wire n_11495;
wire n_1324;
wire n_12034;
wire n_3261;
wire n_12035;
wire n_1544;
wire n_5564;
wire n_12808;
wire n_1327;
wire n_5565;
wire n_414;
wire u15_crac_rd;
wire n_9655;
wire n_5826;
wire n_8436;
wire n_5147;
wire n_8069;
wire n_8472;
wire n_490;
wire oc3_int_set_714;
wire n_10737;
wire n_4477;
wire u8_mem_b2_b_57;
wire n_2138;
wire n_4478;
wire u4_mem_b1_b_83;
wire n_4471;
wire n_2065;
wire n_4476;
wire n_2136;
wire n_4474;
wire n_3872;
wire u8_mem_b3_b_147;
wire n_3869;
wire n_1490;
wire n_3871;
wire u8_mem_b3_b_139;
wire n_4472;
wire n_2207;
wire n_4473;
wire u4_mem_b1_b;
wire n_2116;
wire n_9224;
wire oc0_cfg_970;
wire n_8524;
wire out_slt4;
wire n_10956;
wire n_8606;
wire u13_ints_r_b24_b;
wire n_1245;
wire n_1244;
wire n_12796;
wire u5_mem_b1_b_71;
wire dma_req_o_b2_b;
wire n_982;
wire n_7539;
wire n_2069;
wire n_2068;
wire n_2073;
wire n_2072;
wire n_2070;
wire n_2077;
wire n_2075;
wire n_2074;
wire u9_mem_b3_b_86;
wire n_10701;
wire n_469;
wire n_2218;
wire n_9858;
wire n_3846;
wire n_12166;
wire n_2419;
wire n_1775;
wire n_3549;
wire n_2608;
wire n_675;
wire n_1815;
wire n_581;
wire n_1006;
wire u12_re1;
wire n_2570;
wire n_1209;
wire n_3941;
wire n_2371;
wire n_3942;
wire n_4941;
wire n_2569;
wire n_1224;
wire n_4436;
wire n_9218;
wire n_9290;
wire n_7856;
wire n_7857;
wire n_9221;
wire n_7858;
wire n_9222;
wire n_7859;
wire n_4979;
wire n_7852;
wire n_9214;
wire n_7853;
wire n_9216;
wire n_7854;
wire n_4982;
wire n_7855;
wire n_4444;
wire u4_mem_b1_b_67;
wire n_4977;
wire n_7850;
wire n_4445;
wire n_1940;
wire n_9370;
wire n_2817;
wire n_4625;
wire n_4624;
wire u7_mem_b1_b_83;
wire n_9044;
wire n_9107;
wire n_5487;
wire n_4647;
wire n_5665;
wire u10_mem_b0_b_169;
wire n_5240;
wire u11_mem_b0_b_173;
wire n_5239;
wire n_5251;
wire crac_din_705;
wire n_3983;
wire crac_out_862;
wire n_4681;
wire n_4685;
wire n_4683;
wire oc2_cfg_985;
wire n_4261;
wire n_4686;
wire u13_intm_r_b19_b;
wire u13_ints_r_b19_b;
wire o7_empty;
wire n_7512;
wire n_11658;
wire n_4619;
wire u9_din_tmp_43;
wire n_1448;
wire n_1299;
wire u11_mem_b3_b_78;
wire n_10854;
wire n_8744;
wire n_2976;
wire n_10693;
wire n_1027;
wire n_9236;
wire n_444;
wire n_1383;
wire n_1412;
wire n_1049;
wire n_9687;
wire u8_mem_b3_b_152;
wire n_3768;
wire u4_mem_b0_b_115;
wire n_761;
wire n_11121;
wire o4_we;
wire u3_mem_b3_b_145;
wire n_8368;
wire n_9399;
wire n_1864;
wire n_2723;
wire n_7055;
wire n_5684;
wire n_6158;
wire n_7054;
wire n_5669;
wire n_5801;
wire n_6978;
wire n_5546;
wire n_6981;
wire n_5806;
wire n_7056;
wire n_5700;
wire n_6162;
wire n_7058;
wire n_6164;
wire n_7057;
wire n_5672;
wire n_6979;
wire n_5537;
wire n_5824;
wire n_8894;
wire n_8726;
wire n_8933;
wire n_7053;
wire n_5721;
wire n_5894;
wire u5_mem_b3_b_128;
wire n_9200;
wire n_6556;
wire u11_mem_b3_b_61;
wire n_9274;
wire n_4066;
wire n_10924;
wire u6_mem_b0_b_117;
wire n_8764;
wire n_8908;
wire n_3388;
wire u4_mem_b0_b_93;
wire n_3389;
wire n_2304;
wire n_3391;
wire n_3392;
wire n_1491;
wire u4_mem_b0_b_92;
wire n_9181;
wire n_1547;
wire n_3766;
wire n_11157;
wire n_1325;
wire u5_mem_b3_b_133;
wire n_8810;
wire n_9430;
wire u4_mem_b0_b_99;
wire n_3752;
wire n_7880;
wire u5_mem_b2_b_59;
wire n_7881;
wire u5_mem_b2_b_58;
wire n_8806;
wire u5_mem_b0_b_102;
wire n_3735;
wire n_8807;
wire u5_mem_b0_b_101;
wire n_3737;
wire n_3739;
wire u3_mem_b3_b_143;
wire n_8371;
wire n_9428;
wire n_3734;
wire n_9429;
wire u5_mem_b0_b_103;
wire n_3624;
wire n_7878;
wire n_7879;
wire n_2447;
wire n_8315;
wire u10_mem_b1_b_123;
wire n_10691;
wire n_3929;
wire n_6585;
wire n_2346;
wire u8_mem_b2_b_53;
wire n_12170;
wire u6_mem_b1_b_69;
wire n_8906;
wire u4_wp_b1_b;
wire n_11093;
wire n_8237;
wire u9_mem_b0_b_159;
wire n_10174;
wire n_9148;
wire n_10394;
wire n_9350;
wire n_5096;
wire n_7975;
wire n_7366;
wire n_12303;
wire u9_mem_b2_b_101;
wire n_10283;
wire n_42;
wire ic1_cfg_1035;
wire u9_mem_b1_b_127;
wire n_3908;
wire n_3909;
wire n_3903;
wire n_1564;
wire n_3902;
wire n_3907;
wire n_2269;
wire n_3904;
wire n_2345;
wire n_6014;
wire n_2520;
wire n_2268;
wire n_6465;
wire n_2288;
wire n_4364;
wire u5_mem_b2_b_50;
wire n_2040;
wire n_5007;
wire u6_mem_b1_b_82;
wire n_2650;
wire n_8824;
wire n_5817;
wire n_6201;
wire n_6766;
wire n_6197;
wire n_6195;
wire n_2556;
wire u8_rp_b2_b;
wire u10_mem_b1_b_134;
wire n_1733;
wire n_12304;
wire n_637;
wire o4_empty;
wire n_7513;
wire n_12051;
wire n_2425;
wire n_3080;
wire n_9070;
wire n_4062;
wire n_4063;
wire n_1848;
wire n_4067;
wire u11_din_tmp_47;
wire n_10099;
wire n_1276;
wire n_1816;
wire n_825;
wire n_2420;
wire u10_mem_b3_b_72;
wire n_10225;
wire n_5994;
wire n_6023;
wire n_6630;
wire n_1237;
wire n_6339;
wire n_6575;
wire n_5953;
wire n_5990;
wire n_12061;
wire n_3038;
wire n_4584;
wire u9_din_tmp_46;
wire n_6460;
wire n_1657;
wire n_6428;
wire n_8646;
wire n_8652;
wire n_8651;
wire n_8653;
wire n_8642;
wire u10_mem_b2_b_111;
wire n_10763;
wire n_4848;
wire n_9835;
wire n_9966;
wire n_1549;
wire n_9965;
wire n_9841;
wire n_4850;
wire n_9941;
wire n_9940;
wire n_10875;
wire n_9921;
wire n_9920;
wire n_10876;
wire n_5411;
wire n_10880;
wire n_10372;
wire n_10881;
wire n_10375;
wire n_10879;
wire n_10374;
wire n_5320;
wire n_10378;
wire n_10886;
wire n_10380;
wire n_10885;
wire n_5319;
wire n_10379;
wire n_8390;
wire n_8105;
wire n_8391;
wire n_4517;
wire n_8106;
wire n_11491;
wire n_12607;
wire n_8089;
wire n_9590;
wire n_9487;
wire n_9589;
wire n_9648;
wire n_9549;
wire n_7033;
wire n_1416;
wire n_9876;
wire n_4827;
wire n_9594;
wire n_3994;
wire n_9595;
wire n_2630;
wire n_9592;
wire n_9489;
wire n_10333;
wire n_9844;
wire n_9831;
wire n_9734;
wire n_10777;
wire n_10086;
wire n_8422;
wire n_8091;
wire n_2561;
wire u9_din_tmp_52;
wire u3_mem_b3_b_139;
wire n_90;
wire u10_mem_b1_b_138;
wire n_492;
wire oc0_int_set_708;
wire n_10746;
wire n_5788;
wire u3_mem_b3_b_138;
wire n_11530;
wire n_10163;
wire n_5484;
wire n_10303;
wire n_10162;
wire n_8399;
wire n_8115;
wire n_10169;
wire n_10168;
wire n_10165;
wire n_6863;
wire n_6862;
wire n_5486;
wire n_10167;
wire n_10166;
wire n_6865;
wire n_1477;
wire n_3018;
wire n_3019;
wire n_8907;
wire n_3015;
wire n_3014;
wire n_3016;
wire n_4142;
wire n_11120;
wire n_11463;
wire u8_mem_b0_b_94;
wire u11_din_tmp_50;
wire n_10096;
wire n_7523;
wire u3_mem_b2_b_32;
wire n_8396;
wire oc4_cfg_1005;
wire n_9283;
wire n_8281;
wire u5_rp_b2_b;
wire n_1719;
wire n_6859;
wire n_6879;
wire u11_mem_b0_b_180;
wire u11_mem_b1_b_121;
wire n_10552;
wire u9_mem_b3_b_78;
wire n_10709;
wire n_11661;
wire n_12272;
wire n_3493;
wire n_12091;
wire n_3495;
wire n_3497;
wire n_4243;
wire n_9273;
wire n_1247;
wire n_1246;
wire n_1415;
wire n_4240;
wire u7_mem_b1_b_82;
wire u9_mem_b1_b_130;
wire n_10397;
wire n_11002;
wire n_11163;
wire n_11512;
wire n_11513;
wire n_10968;
wire n_11153;
wire n_10969;
wire n_11160;
wire n_11508;
wire n_11509;
wire n_11161;
wire n_11510;
wire n_11511;
wire n_11150;
wire n_10986;
wire n_11151;
wire n_10993;
wire n_5372;
wire u9_mem_b3_b_79;
wire n_9246;
wire n_12214;
wire n_9633;
wire n_9737;
wire n_11699;
wire n_2833;
wire n_4454;
wire n_1962;
wire n_5117;
wire u7_mem_b1_b_63;
wire n_2738;
wire n_4459;
wire n_2063;
wire n_2208;
wire n_4461;
wire u4_mem_b1_b_60;
wire n_2184;
wire n_4455;
wire n_4456;
wire n_4458;
wire u4_mem_b1_b_81;
wire n_2061;
wire n_3209;
wire u5_mem_b3_b_139;
wire u11_mem_b0_b_167;
wire n_10899;
wire n_1562;
wire u9_mem_b0_b_172;
wire n_2529;
wire n_6612;
wire n_11023;
wire u9_mem_b2_b_115;
wire i3_dout_565;
wire n_4046;
wire n_232;
wire n_8320;
wire n_4453;
wire n_8031;
wire n_8033;
wire n_8321;
wire n_8325;
wire n_8035;
wire n_8324;
wire n_8034;
wire n_8327;
wire n_8037;
wire n_8326;
wire n_8036;
wire n_9347;
wire n_8317;
wire n_8029;
wire n_9058;
wire n_12527;
wire n_12526;
wire n_12528;
wire n_12529;
wire n_283;
wire u5_mem_b1_b;
wire n_9317;
wire n_2469;
wire n_4854;
wire n_4266;
wire n_754;
wire n_3560;
wire n_923;
wire n_5645;
wire n_4153;
wire n_4640;
wire n_3561;
wire n_10160;
wire n_9235;
wire n_7871;
wire n_9237;
wire n_7872;
wire n_4353;
wire n_9264;
wire n_7875;
wire n_9241;
wire n_4354;
wire n_7876;
wire n_4351;
wire n_7873;
wire n_4352;
wire n_7874;
wire n_9244;
wire n_4355;
wire n_9245;
wire n_4356;
wire n_9242;
wire n_4308;
wire n_7877;
wire n_9243;
wire n_3467;
wire n_4073;
wire n_10781;
wire n_10903;
wire n_10973;
wire n_10573;
wire n_10974;
wire n_10977;
wire n_10587;
wire n_10979;
wire n_10589;
wire n_9962;
wire n_12656;
wire n_1457;
wire n_9492;
wire n_2649;
wire i6_dout_645;
wire n_4019;
wire n_4735;
wire n_10402;
wire n_3470;
wire rf_we;
wire n_6041;
wire n_5288;
wire n_5283;
wire u10_mem_b2_b_110;
wire n_4742;
wire n_5281;
wire n_5280;
wire n_4741;
wire oc5_cfg_1015;
wire n_5279;
wire u13_intm_r_b10_b;
wire crac_din_701;
wire u8_mem_b0_b_104;
wire n_748;
wire n_3469;
wire u3_mem_b1_b_78;
wire n_11752;
wire u2_bit_clk_r;
wire n_9773;
wire n_11134;
wire n_4821;
wire u9_mem_b1_b_135;
wire n_10304;
wire n_1196;
wire n_9346;
wire n_6896;
wire n_6908;
wire n_6003;
wire n_6577;
wire n_6576;
wire n_1667;
wire n_6426;
wire n_1005;
wire n_8899;
wire n_6739;
wire n_121;
wire n_6876;
wire u9_mem_b1_b_122;
wire oc4_int_set;
wire n_9848;
wire u10_din_tmp_48;
wire n_9865;
wire n_12850;
wire n_3538;
wire n_2983;
wire n_1669;
wire n_1668;
wire n_6966;
wire n_5784;
wire n_6965;
wire n_5783;
wire n_6964;
wire oc0_cfg_969;
wire n_5782;
wire n_6963;
wire n_5781;
wire n_6962;
wire n_5780;
wire n_6961;
wire oc1_cfg_974;
wire n_5779;
wire n_6960;
wire n_5761;
wire n_6959;
wire n_5786;
wire n_6958;
wire n_5777;
wire n_6038;
wire n_6037;
wire u10_mem_b1_b_133;
wire n_3383;
wire u3_mem_b2_b_31;
wire n_3381;
wire n_2238;
wire u13_ints_r_b8_b;
wire n_11011;
wire n_8277;
wire n_1977;
wire n_1466;
wire n_2239;
wire n_2925;
wire n_7652;
wire n_7653;
wire n_7654;
wire n_7646;
wire n_7647;
wire n_7648;
wire u7_mem_b3_b_134;
wire n_7649;
wire u7_mem_b3_b_138;
wire n_7645;
wire n_10278;
wire u10_mem_b0_b_164;
wire u10_din_tmp_49;
wire n_9863;
wire out_slt_25;
wire n_1031;
wire i6_dout_652;
wire n_7860;
wire n_7861;
wire n_7862;
wire n_7863;
wire n_7864;
wire n_7865;
wire n_7866;
wire u9_wp_b1_b;
wire u10_mem_b2_b;
wire n_665;
wire oc2_int_set_711;
wire u8_mem_b2_b_43;
wire n_12262;
wire n_12269;
wire u3_mem_b2_b_39;
wire n_753;
wire u11_mem_b0_b;
wire n_10821;
wire n_1395;
wire n_10670;
wire u9_mem_b2_b_112;
wire n_2397;
wire u3_mem_b3_b_132;
wire n_2945;
wire u7_mem_b2_b_31;
wire n_11052;
wire n_4029;
wire u13_intm_r_b4_b;
wire n_8492;
wire u9_mem_b0_b_155;
wire u10_mem_b3_b_71;
wire u10_mem_b2_b_101;
wire n_36;
wire n_10253;
wire n_3938;
wire n_4220;
wire n_4626;
wire n_2354;
wire n_3081;
wire n_3937;
wire u9_mem_b0_b_156;
wire n_10143;
wire n_6916;
wire n_3373;
wire n_1925;
wire n_6952;
wire n_2259;
wire n_6771;
wire n_6206;
wire n_6210;
wire n_6209;
wire n_5594;
wire n_11597;
wire n_6772;
wire n_6774;
wire n_6763;
wire n_1014;
wire n_6208;
wire n_6207;
wire n_431;
wire n_9083;
wire n_8982;
wire u10_mem_b1_b_122;
wire u9_mem_b3_b_80;
wire n_6424;
wire u11_mem_b3_b_69;
wire n_6633;
wire u10_mem_b2_b_90;
wire u9_mem_b3_b_66;
wire u9_mem_b3_b_68;
wire n_403;
wire u3_mem_b2_b_38;
wire n_808;
wire n_11180;
wire n_8296;
wire n_603;
wire n_5;
wire n_696;
wire n_463;
wire n_1054;
wire n_1367;
wire n_10678;
wire n_5419;
wire n_9993;
wire n_5428;
wire n_10393;
wire n_9081;
wire u9_mem_b2_b_111;
wire n_10690;
wire n_5515;
wire n_10688;
wire n_5513;
wire n_10686;
wire n_5360;
wire n_10004;
wire n_10685;
wire n_5358;
wire n_10684;
wire n_5353;
wire n_10002;
wire n_5511;
wire n_10001;
wire n_5507;
wire n_10000;
wire n_10680;
wire n_5505;
wire n_9999;
wire n_9449;
wire n_1444;
wire n_10449;
wire n_6044;
wire n_590;
wire n_929;
wire n_1038;
wire n_10145;
wire n_6850;
wire n_6848;
wire n_6847;
wire n_6395;
wire n_10141;
wire n_6846;
wire n_10148;
wire n_6858;
wire n_6857;
wire n_10147;
wire n_6855;
wire n_10822;
wire n_9907;
wire n_10146;
wire n_6853;
wire n_10140;
wire n_9843;
wire n_10139;
wire n_8874;
wire n_4861;
wire n_7947;
wire n_8329;
wire n_8041;
wire n_7751;
wire n_7088;
wire n_9121;
wire n_8876;
wire n_8076;
wire n_2049;
wire n_7753;
wire u6_mem_b3_b_136;
wire u6_rp_b0_b;
wire n_11113;
wire n_5916;
wire n_8717;
wire n_8154;
wire n_7571;
wire n_1134;
wire n_8869;
wire n_4291;
wire n_7616;
wire n_1063;
wire n_9088;
wire n_4417;
wire n_7995;
wire n_6300;
wire n_5694;
wire u5_wp_b2_b;
wire n_9467;
wire n_10134;
wire n_8165;
wire u8_mem_b3_b_132;
wire n_8275;
wire n_4418;
wire n_7996;
wire u6_mem_b1_b_66;
wire n_9152;
wire n_9025;
wire n_8270;
wire n_4411;
wire n_7991;
wire u11_mem_b1_b_134;
wire n_10842;
wire n_4410;
wire n_7990;
wire n_9698;
wire n_9523;
wire n_9767;
wire n_9600;
wire n_9658;
wire n_9700;
wire n_9524;
wire n_9613;
wire n_7275;
wire n_6129;
wire n_10089;
wire n_9504;
wire n_9755;
wire u15_rdd2;
wire n_9883;
wire n_7325;
wire n_6833;
wire n_6126;
wire n_9847;
wire n_9696;
wire n_9522;
wire n_9652;
wire n_3511;
wire n_7320;
wire n_11539;
wire n_11540;
wire n_10400;
wire n_9561;
wire n_9837;
wire n_6807;
wire n_6078;
wire n_1695;
wire n_6080;
wire n_4195;
wire n_3108;
wire n_2277;
wire n_4259;
wire n_4144;
wire n_2972;
wire n_2260;
wire n_4252;
wire n_4147;
wire n_3393;
wire n_2348;
wire n_4260;
wire n_6081;
wire n_9029;
wire n_7424;
wire n_8372;
wire n_8369;
wire n_4852;
wire n_10538;
wire n_3945;
wire n_12270;
wire n_1294;
wire n_12278;
wire n_2504;
wire n_5957;
wire u9_mem_b1_b_132;
wire n_10307;
wire n_5194;
wire n_2432;
wire n_3315;
wire n_6263;
wire n_6165;
wire n_4098;
wire u11_din_tmp_56;
wire n_10245;
wire n_10778;
wire u9_mem_b3_b_69;
wire n_10258;
wire n_8352;
wire n_7834;
wire n_7592;
wire n_8350;
wire n_8147;
wire n_8349;
wire n_4485;
wire n_7558;
wire n_8348;
wire n_4960;
wire n_4855;
wire n_7559;
wire n_4345;
wire n_8066;
wire n_8345;
wire n_8056;
wire n_8344;
wire n_4381;
wire n_8055;
wire n_8343;
wire n_4138;
wire n_4111;
wire n_5241;
wire n_4237;
wire n_5242;
wire n_4205;
wire n_3949;
wire n_4643;
wire n_3950;
wire n_4645;
wire n_4644;
wire n_4642;
wire n_2994;
wire n_5238;
wire n_4202;
wire n_4368;
wire n_7893;
wire n_9262;
wire n_4276;
wire n_7894;
wire n_4369;
wire n_7895;
wire n_9265;
wire n_4371;
wire n_7896;
wire n_9266;
wire n_4372;
wire n_7897;
wire n_9267;
wire n_4373;
wire n_7898;
wire n_9268;
wire n_4374;
wire n_7899;
wire n_4542;
wire n_7900;
wire n_12827;
wire n_2246;
wire n_3539;
wire n_5678;
wire n_6144;
wire n_3375;
wire n_3119;
wire n_1508;
wire n_5677;
wire n_5803;
wire n_11467;
wire n_11468;
wire n_2245;
wire n_2395;
wire n_5536;
wire n_9258;
wire n_4365;
wire n_7891;
wire n_9259;
wire n_4367;
wire n_7892;
wire n_12817;
wire n_4722;
wire u13_intm_r_b22_b;
wire n_8374;
wire n_5132;
wire n_8090;
wire n_4723;
wire n_3989;
wire n_5197;
wire n_4143;
wire n_3041;
wire u13_intm_r_b24_b;
wire n_4311;
wire u7_mem_b2_b_54;
wire n_4720;
wire n_7969;
wire u11_din_tmp_54;
wire n_6372;
wire n_5274;
wire u13_intm_r_b25_b;
wire n_4303;
wire n_2019;
wire n_5093;
wire n_8087;
wire n_5634;
wire n_4102;
wire n_2606;
wire n_7964;
wire n_8370;
wire n_5131;
wire n_8061;
wire n_8366;
wire n_5123;
wire n_7967;
wire n_8554;
wire n_1216;
wire n_5759;
wire n_5171;
wire n_4580;
wire n_8290;
wire n_6106;
wire n_5461;
wire n_5205;
wire n_6105;
wire n_4610;
wire n_6104;
wire n_12060;
wire n_5168;
wire n_9457;
wire n_5758;
wire n_4574;
wire n_5172;
wire n_12513;
wire n_12514;
wire n_12506;
wire n_12507;
wire n_12508;
wire u4_mem_b3_b_146;
wire n_9337;
wire n_12509;
wire n_9768;
wire n_9660;
wire n_9699;
wire n_9612;
wire n_7519;
wire n_9702;
wire n_9701;
wire n_9615;
wire n_11672;
wire n_11673;
wire n_9473;
wire n_10403;
wire n_9657;
wire n_9646;
wire n_9697;
wire n_9588;
wire n_1388;
wire n_996;
wire n_6536;
wire n_6535;
wire n_6880;
wire n_6877;
wire n_6529;
wire n_2819;
wire n_2832;
wire u11_mem_b0_b_176;
wire u11_mem_b2_b_111;
wire u14_n_133;
wire n_12459;
wire n_7796;
wire n_6046;
wire n_5671;
wire n_6234;
wire n_6990;
wire n_5547;
wire n_6989;
wire n_5555;
wire n_5856;
wire n_7092;
wire n_5838;
wire n_6991;
wire n_5548;
wire n_5836;
wire n_7090;
wire n_6215;
wire n_5692;
wire n_6212;
wire n_7183;
wire n_7091;
wire n_5693;
wire n_6217;
wire n_7267;
wire n_6733;
wire n_5614;
wire u10_mem_b2_b_115;
wire n_10446;
wire n_7666;
wire n_7669;
wire n_7670;
wire n_7667;
wire n_7668;
wire n_7451;
wire n_7674;
wire n_7671;
wire n_7672;
wire n_8365;
wire u8_mem_b1_b_64;
wire n_4212;
wire n_4214;
wire u7_mem_b1_b_85;
wire n_3358;
wire n_1364;
wire n_3353;
wire n_9002;
wire u10_mem_b3_b_82;
wire n_7919;
wire n_7920;
wire u5_mem_b1_b_85;
wire n_4880;
wire n_7929;
wire n_7930;
wire n_7925;
wire u5_mem_b1_b_80;
wire n_7923;
wire u5_mem_b1_b_82;
wire n_7924;
wire n_7921;
wire u5_mem_b1_b_84;
wire n_7922;
wire u5_mem_b1_b_83;
wire n_8389;
wire n_4859;
wire n_8104;
wire i3_dout_590;
wire n_4049;
wire n_12464;
wire n_12454;
wire n_12460;
wire n_10298;
wire n_9172;
wire n_2255;
wire n_8854;
wire n_503;
wire n_1861;
wire u6_mem_b3_b_130;
wire n_8401;
wire u10_mem_b3_b_57;
wire n_10223;
wire n_12612;
wire u3_mem_b0_b_102;
wire u9_mem_b2_b_118;
wire n_12613;
wire n_10212;
wire n_4020;
wire n_2932;
wire n_8382;
wire n_4955;
wire n_8096;
wire n_11656;
wire n_3248;
wire n_3547;
wire n_9310;
wire n_5510;
wire n_1690;
wire u3_rp_b0_b;
wire n_12834;
wire n_2814;
wire u4_mem_b2_b_32;
wire n_2192;
wire n_2182;
wire n_2815;
wire n_2190;
wire n_2196;
wire n_2816;
wire n_2195;
wire n_11503;
wire u10_mem_b3_b_62;
wire n_4089;
wire n_10408;
wire n_9555;
wire n_4023;
wire u4_mem_b0_b_91;
wire n_8829;
wire n_10893;
wire u10_mem_b0_b_172;
wire n_10129;
wire n_6048;
wire n_11164;
wire u10_mem_b1_b_121;
wire u8_mem_b2_b_50;
wire n_9132;
wire u9_mem_b0_b_160;
wire n_2509;
wire n_3599;
wire n_694;
wire u13_ints_r_b10_b;
wire n_450;
wire n_914;
wire n_10850;
wire n_5501;
wire n_10350;
wire n_5503;
wire n_5497;
wire n_10352;
wire n_10851;
wire n_5493;
wire n_10351;
wire n_10846;
wire n_5509;
wire n_10346;
wire n_10845;
wire n_5523;
wire n_10345;
wire n_10848;
wire n_5499;
wire n_10348;
wire n_5525;
wire n_10347;
wire n_9974;
wire n_10661;
wire n_9973;
wire n_6598;
wire u10_mem_b3_b_67;
wire n_8445;
wire n_4702;
wire n_1035;
wire n_1908;
wire n_9567;
wire n_9448;
wire n_9447;
wire n_729;
wire n_2896;
wire n_3611;
wire n_10447;
wire n_10131;
wire n_5956;
wire n_10448;
wire n_5954;
wire n_6361;
wire n_10132;
wire n_5958;
wire n_10814;
wire n_6364;
wire n_9640;
wire u10_mem_b2_b_89;
wire n_8938;
wire n_11650;
wire n_792;
wire u13_intm_r_b1_b;
wire u8_mem_b1_b;
wire n_1462;
wire u8_mem_b3_b_146;
wire n_693;
wire i3_dout_591;
wire n_4048;
wire u11_mem_b2_b_103;
wire n_5966;
wire n_2574;
wire n_838;
wire u9_mem_b2_b_98;
wire u10_mem_b1_b_120;
wire u11_mem_b2_b;
wire u11_mem_b3_b_86;
wire n_12539;
wire n_12537;
wire n_12538;
wire n_12533;
wire n_5723;
wire n_6134;
wire n_6131;
wire u13_intm_r_b27_b;
wire u13_intm_r_b28_b;
wire u4_mem_b0_b_94;
wire n_2893;
wire u11_mem_b3_b_62;
wire n_10828;
wire u6_mem_b2_b_56;
wire n_3686;
wire n_10943;
wire n_7264;
wire n_5932;
wire n_6121;
wire n_7127;
wire n_5933;
wire n_5768;
wire n_7128;
wire n_5934;
wire n_5769;
wire n_7265;
wire n_6314;
wire n_6092;
wire n_7318;
wire n_6130;
wire n_7266;
wire n_5773;
wire n_7132;
wire n_5774;
wire n_7129;
wire n_5935;
wire n_5770;
wire n_7130;
wire n_5936;
wire n_5771;
wire n_5722;
wire n_11646;
wire n_11647;
wire n_3166;
wire n_3532;
wire u13_intm_r_b18_b;
wire n_3925;
wire n_1248;
wire n_5389;
wire n_1687;
wire n_3923;
wire n_4038;
wire n_1572;
wire n_1571;
wire n_5388;
wire n_5387;
wire n_6157;
wire n_12004;
wire n_12005;
wire n_3336;
wire n_2450;
wire n_2559;
wire n_3919;
wire n_9031;
wire n_730;
wire u11_mem_b3_b_70;
wire n_10457;
wire n_8502;
wire n_664;
wire n_4816;
wire ic0_int_set;
wire n_7480;
wire oc5_int_set;
wire n_3277;
wire u7_mem_b2_b_30;
wire n_9420;
wire n_2372;
wire n_8268;
wire n_4409;
wire n_7989;
wire n_8153;
wire u4_mem_b2_b_35;
wire n_8162;
wire n_7997;
wire n_8157;
wire u8_mem_b3_b_138;
wire n_8156;
wire n_4414;
wire n_7993;
wire n_1319;
wire n_886;
wire n_8474;
wire n_4651;
wire n_5467;
wire n_1894;
wire n_5466;
wire n_5244;
wire n_4650;
wire n_5304;
wire n_4649;
wire n_5243;
wire n_4193;
wire n_4648;
wire n_3061;
wire n_3953;
wire n_1021;
wire n_635;
wire n_2989;
wire n_9294;
wire n_5027;
wire n_9296;
wire n_5028;
wire n_5025;
wire n_9293;
wire n_5026;
wire n_7917;
wire n_5024;
wire n_7918;
wire n_9285;
wire n_7915;
wire n_7916;
wire n_7913;
wire n_7914;
wire n_725;
wire u13_intm_r_b11_b;
wire u13_intm_r_b12_b;
wire n_8394;
wire n_8245;
wire u11_mem_b0_b_163;
wire n_2066;
wire n_8952;
wire u13_ints_r_b25_b;
wire u13_ints_r_b26_b;
wire n_8655;
wire n_4297;
wire u4_mem_b1_b_65;
wire n_2481;
wire n_4875;
wire n_2890;
wire n_4299;
wire n_4876;
wire n_4877;
wire n_3446;
wire n_4878;
wire n_3444;
wire n_4879;
wire n_4300;
wire n_2177;
wire n_8511;
wire n_8519;
wire n_8512;
wire n_8517;
wire n_8518;
wire n_8520;
wire n_8514;
wire n_3997;
wire n_2498;
wire n_3346;
wire n_4978;
wire n_3123;
wire u11_mem_b2_b_88;
wire u9_din_tmp_53;
wire i4_dout_598;
wire u9_din_tmp_54;
wire n_6758;
wire n_3809;
wire n_1709;
wire n_3812;
wire n_5764;
wire n_4587;
wire n_5183;
wire n_5584;
wire n_3967;
wire n_6119;
wire n_5458;
wire n_6117;
wire n_5557;
wire n_5765;
wire n_5254;
wire n_3978;
wire n_5538;
wire n_5767;
wire n_5167;
wire n_5166;
wire n_6122;
wire n_5214;
wire n_5460;
wire n_2098;
wire n_3029;
wire crac_din_692;
wire n_1202;
wire n_11008;
wire n_10775;
wire n_10806;
wire n_9616;
wire n_5840;
wire n_5832;
wire n_9659;
wire n_5828;
wire n_9656;
wire n_8845;
wire n_1153;
wire n_667;
wire n_11612;
wire n_8636;
wire n_2270;
wire n_6626;
wire n_6634;
wire n_6934;
wire n_6933;
wire n_6636;
wire n_6635;
wire n_6936;
wire n_6935;
wire n_6631;
wire n_6932;
wire n_6931;
wire n_12354;
wire n_11843;
wire n_2827;
wire n_6753;
wire n_10110;
wire n_10339;
wire n_1103;
wire n_7687;
wire n_7688;
wire n_7689;
wire u7_mem_b1_b_64;
wire n_7690;
wire n_7691;
wire n_7692;
wire u7_mem_b1_b_89;
wire n_7693;
wire u3_mem_b1_b_83;
wire n_7685;
wire oc3_cfg;
wire u7_mem_b0_b_94;
wire n_9392;
wire n_8253;
wire n_9037;
wire n_9470;
wire out_slt_24;
wire n_6987;
wire n_7080;
wire n_8671;
wire n_9480;
wire n_11841;
wire n_7177;
wire n_6084;
wire n_4208;
wire n_8670;
wire n_7542;
wire n_5675;
wire n_5816;
wire n_7256;
wire n_7904;
wire n_7906;
wire u5_mem_b1_b_68;
wire n_7908;
wire u5_mem_b1_b_67;
wire n_7901;
wire n_7902;
wire n_7903;
wire n_10136;
wire n_4056;
wire n_9232;
wire n_3806;
wire u7_mem_b0_b_101;
wire n_11122;
wire n_5447;
wire n_7341;
wire n_7343;
wire n_7342;
wire n_1133;
wire n_7027;
wire n_7019;
wire n_7022;
wire n_5623;
wire n_8795;
wire n_9681;
wire n_6740;
wire n_5868;
wire u6_mem_b2_b_30;
wire n_9122;
wire u7_mem_b1_b_80;
wire n_9047;
wire n_11072;
wire n_9199;
wire n_10127;
wire n_2203;
wire n_2205;
wire u8_mem_b0_b_120;
wire n_9375;
wire n_2822;
wire n_2823;
wire n_421;
wire n_6742;
wire u10_mem_b2_b_100;
wire u9_mem_b0_b_168;
wire u8_mem_b1_b_67;
wire n_11129;
wire oc4_cfg_1009;
wire n_1126;
wire n_9104;
wire u5_mem_b2_b_54;
wire n_9253;
wire u9_mem_b1_b_144;
wire n_4752;
wire n_5489;
wire n_5488;
wire n_4654;
wire n_5346;
wire n_5345;
wire n_5344;
wire n_5348;
wire n_5340;
wire n_5339;
wire n_4748;
wire u9_mem_b2_b_108;
wire n_1845;
wire n_12172;
wire n_5582;
wire u7_rp_b1_b;
wire n_11085;
wire n_6744;
wire n_9023;
wire n_8875;
wire n_1163;
wire n_4766;
wire n_9980;
wire n_10667;
wire n_9979;
wire n_10672;
wire n_5291;
wire n_9984;
wire n_5289;
wire n_9983;
wire n_9982;
wire n_10669;
wire n_5356;
wire n_9981;
wire n_5297;
wire n_10360;
wire n_5496;
wire n_10859;
wire n_5301;
wire n_10359;
wire n_10673;
wire n_4746;
wire n_9985;
wire n_8024;
wire n_5617;
wire n_7686;
wire u7_mem_b1_b_67;
wire u5_mem_b2_b_34;
wire n_1146;
wire n_1007;
wire n_1309;
wire n_8664;
wire n_1023;
wire n_9511;
wire n_8669;
wire n_1302;
wire n_9510;
wire n_8666;
wire n_1373;
wire n_9512;
wire n_1375;
wire n_9513;
wire u14_u7_en_out_l2;
wire n_8364;
wire u11_mem_b2_b_90;
wire n_8465;
wire n_7838;
wire u4_mem_b1_b_86;
wire n_7311;
wire n_6820;
wire n_11031;
wire n_11621;
wire n_11622;
wire n_1809;
wire u7_mem_b0_b_97;
wire n_8455;
wire n_7618;
wire n_8028;
wire n_11028;
wire n_11731;
wire n_11732;
wire n_3845;
wire n_6789;
wire n_6791;
wire n_7248;
wire n_6223;
wire n_6238;
wire n_6236;
wire n_6235;
wire n_6786;
wire n_8693;
wire u11_mem_b1_b_128;
wire n_10731;
wire n_9226;
wire n_3078;
wire n_6111;
wire n_6112;
wire n_11019;
wire n_11637;
wire n_11638;
wire n_11992;
wire n_11993;
wire n_6116;
wire n_11022;
wire n_12016;
wire n_12017;
wire n_11629;
wire n_11024;
wire n_11735;
wire n_11026;
wire n_11625;
wire n_11027;
wire n_11733;
wire n_11734;
wire n_3360;
wire oc3_cfg_1000;
wire n_9435;
wire n_3550;
wire i6_dout_632;
wire n_4003;
wire u11_mem_b2_b_91;
wire n_10498;
wire u10_mem_b2_b_114;
wire u4_rp_b1_b;
wire n_2257;
wire n_2995;
wire n_4256;
wire n_2997;
wire n_2996;
wire u3_mem_b2_b_44;
wire n_2634;
wire u3_mem_b1_b_68;
wire n_4050;
wire n_1705;
wire n_1729;
wire n_1726;
wire n_4052;
wire n_1563;
wire n_1735;
wire n_1734;
wire n_1718;
wire n_4045;
wire n_2508;
wire n_1858;
wire n_1725;
wire n_1722;
wire n_4047;
wire n_2501;
wire n_1720;
wire n_2117;
wire n_4044;
wire n_1717;
wire n_2505;
wire n_4043;
wire n_1714;
wire n_1712;
wire n_2185;
wire n_11084;
wire n_9859;
wire n_4209;
wire n_3344;
wire n_1475;
wire n_2341;
wire n_7076;
wire n_5685;
wire n_6193;
wire n_478;
wire n_11443;
wire n_10758;
wire n_741;
wire n_7531;
wire n_872;
wire n_4706;
wire n_5385;
wire n_12334;
wire n_11507;
wire n_8295;
wire n_7713;
wire n_8293;
wire n_4432;
wire n_8016;
wire n_9062;
wire n_7718;
wire n_7717;
wire n_2316;
wire n_8132;
wire n_8131;
wire n_7707;
wire n_9048;
wire n_7706;
wire u11_mem_b3_b_81;
wire n_10920;
wire n_2888;
wire n_8592;
wire n_5542;
wire n_5541;
wire u8_mem_b2_b_30;
wire n_2002;
wire n_5687;
wire n_4196;
wire n_6228;
wire n_2289;
wire n_1531;
wire n_4210;
wire n_1275;
wire n_1533;
wire n_6072;
wire n_5245;
wire n_4238;
wire n_9884;
wire n_9312;
wire n_5042;
wire n_7936;
wire n_9313;
wire n_5043;
wire n_7938;
wire n_4384;
wire n_5064;
wire n_7950;
wire n_9320;
wire n_7951;
wire n_9321;
wire n_5067;
wire n_9314;
wire n_5023;
wire n_7939;
wire n_5046;
wire n_7941;
wire n_9316;
wire n_5047;
wire n_7942;
wire n_5049;
wire n_7943;
wire n_1502;
wire n_12479;
wire n_12482;
wire n_8392;
wire n_3963;
wire n_4283;
wire n_4284;
wire n_2122;
wire n_1686;
wire n_1683;
wire n_4290;
wire n_1987;
wire u8_mem_b2_b_48;
wire n_2176;
wire n_1556;
wire n_4289;
wire n_1936;
wire n_2119;
wire n_4285;
wire n_2202;
wire n_4286;
wire n_1960;
wire n_2043;
wire n_3483;
wire u7_mem_b0_b_110;
wire n_12499;
wire n_12500;
wire n_9947;
wire n_6808;
wire n_6806;
wire n_6804;
wire n_6801;
wire n_9752;
wire n_1435;
wire u11_mem_b2_b_116;
wire n_10862;
wire n_2363;
wire u7_mem_b0_b_107;
wire n_8747;
wire n_2580;
wire n_2579;
wire n_6250;
wire n_7441;
wire n_630;
wire n_6124;
wire n_6282;
wire n_5909;
wire n_5811;
wire n_6590;
wire n_6588;
wire n_6278;
wire n_6280;
wire u9_mem_b0_b_167;
wire n_10765;
wire n_8957;
wire n_2417;
wire n_831;
wire n_2418;
wire n_2423;
wire n_2424;
wire n_8763;
wire n_8912;
wire n_2416;
wire u6_mem_b3_b_122;
wire n_6600;
wire n_6917;
wire n_6915;
wire n_6597;
wire n_6595;
wire n_9179;
wire n_4382;
wire n_2214;
wire n_1663;
wire n_162;
wire n_5504;
wire o8_we;
wire n_7024;
wire n_6511;
wire n_3527;
wire n_2532;
wire n_1661;
wire n_6507;
wire n_6421;
wire n_2533;
wire n_11165;
wire u4_mem_b1_b_64;
wire n_8308;
wire n_9050;
wire u11_mem_b2_b_108;
wire n_10873;
wire n_7716;
wire n_7715;
wire n_7710;
wire n_7708;
wire n_7705;
wire n_7435;
wire n_7436;
wire n_9617;
wire n_11613;
wire n_7122;
wire n_7065;
wire n_3333;
wire n_12038;
wire u8_mem_b2_b_31;
wire n_3338;
wire n_4206;
wire n_12036;
wire u8_mem_b2_b_44;
wire n_5317;
wire n_2336;
wire u10_mem_b1_b_119;
wire n_8739;
wire n_9396;
wire u7_mem_b0_b_112;
wire n_3641;
wire u10_din_tmp_56;
wire n_9854;
wire n_8745;
wire u7_mem_b0_b_108;
wire n_3564;
wire n_3644;
wire n_3645;
wire n_8740;
wire u7_mem_b0_b_111;
wire n_3568;
wire n_8742;
wire n_3642;
wire n_3566;
wire n_9398;
wire n_2635;
wire n_10173;
wire n_9065;
wire n_7376;
wire u11_mem_b1_b_145;
wire n_1192;
wire crac_din_704;
wire n_7389;
wire n_7357;
wire n_7388;
wire in_valid_s_b2_b;
wire n_11038;
wire n_11155;
wire n_3198;
wire n_4167;
wire n_1074;
wire crac_din;
wire n_4809;
wire n_1612;
wire n_525;
wire n_12667;
wire n_11923;
wire n_4016;
wire n_1621;
wire n_1617;
wire n_10226;
wire n_3092;
wire n_2796;
wire o6_empty;
wire n_7438;
wire n_2791;
wire u3_mem_b3_b_137;
wire n_2162;
wire n_2161;
wire n_4951;
wire n_2694;
wire n_4343;
wire n_2084;
wire u3_mem_b3_b_135;
wire n_3478;
wire u9_mem_b2_b_91;
wire n_10270;
wire n_3091;
wire u11_din_tmp_42;
wire n_10105;
wire n_3090;
wire n_5763;
wire n_3957;
wire n_10730;
wire n_4658;
wire n_6062;
wire n_4655;
wire n_5351;
wire n_5350;
wire n_5500;
wire n_4652;
wire n_256;
wire n_2307;
wire n_337;
wire n_3927;
wire n_1689;
wire n_1691;
wire n_314;
wire n_10057;
wire n_600;
wire n_9882;
wire n_7260;
wire n_7096;
wire n_7258;
wire n_7116;
wire n_7262;
wire n_7047;
wire n_7126;
wire n_7099;
wire n_9803;
wire n_9710;
wire n_12008;
wire n_7279;
wire n_7105;
wire n_2303;
wire n_3185;
wire n_3184;
wire u3_mem_b2_b_56;
wire n_3186;
wire n_703;
wire n_10362;
wire n_10361;
wire n_9986;
wire n_87;
wire n_5013;
wire n_2758;
wire n_5929;
wire n_10668;
wire n_1042;
wire n_6891;
wire n_11667;
wire oc4_cfg_1006;
wire n_8280;
wire u6_mem_b1_b_72;
wire u10_mem_b0_b_159;
wire n_8917;
wire n_4870;
wire n_7600;
wire n_1570;
wire n_7949;
wire n_4281;
wire n_7602;
wire n_10708;
wire n_4869;
wire n_7597;
wire n_8910;
wire n_7564;
wire n_4280;
wire n_7599;
wire n_5800;
wire n_8914;
wire n_7598;
wire n_334;
wire n_4868;
wire n_6298;
wire n_9348;
wire n_5095;
wire n_4279;
wire n_7124;
wire n_7244;
wire n_6145;
wire n_6283;
wire n_7245;
wire n_7246;
wire n_6297;
wire u9_mem_b0_b_151;
wire n_10152;
wire n_2471;
wire n_9082;
wire n_9080;
wire n_9078;
wire n_5101;
wire n_7732;
wire n_6919;
wire u11_mem_b0_b_179;
wire n_8151;
wire n_8266;
wire n_5580;
wire u11_mem_b3_b_74;
wire n_7983;
wire u4_mem_b1_b_69;
wire n_3010;
wire n_8150;
wire u8_mem_b3_b_144;
wire n_7338;
wire n_5276;
wire n_2886;
wire n_4761;
wire u10_mem_b0_b_168;
wire n_10677;
wire n_8260;
wire n_7980;
wire n_7981;
wire n_10417;
wire u7_mem_b2_b_57;
wire u14_u6_full_empty_r;
wire n_12799;
wire n_12800;
wire n_1338;
wire n_4822;
wire n_2554;
wire n_5727;
wire n_8259;
wire n_5099;
wire n_7979;
wire n_4823;
wire n_1840;
wire n_2555;
wire n_11662;
wire n_11663;
wire n_3533;
wire n_3431;
wire n_7524;
wire n_1624;
wire n_4027;
wire n_11049;
wire n_9301;
wire n_3999;
wire n_6809;
wire n_5188;
wire n_10554;
wire n_5187;
wire n_1811;
wire n_3840;
wire n_6694;
wire n_2871;
wire n_2984;
wire i3_dout_567;
wire n_4033;
wire n_2464;
wire n_3122;
wire n_10157;
wire n_5186;
wire n_3004;
wire n_9033;
wire n_4893;
wire n_5009;
wire n_4892;
wire n_9028;
wire n_9026;
wire n_5070;
wire n_8112;
wire n_8110;
wire n_8114;
wire n_8113;
wire n_8116;
wire n_8118;
wire n_8117;
wire n_8120;
wire u3_mem_b2_b_55;
wire n_8119;
wire n_5897;
wire n_5805;
wire n_4487;
wire n_2165;
wire n_5895;
wire n_4486;
wire u3_mem_b2_b_46;
wire n_3032;
wire n_3877;
wire u8_mem_b3_b_130;
wire n_1470;
wire n_9772;
wire n_7012;
wire n_6403;
wire n_4659;
wire n_10756;
wire u8_mem_b0_b_107;
wire n_9381;
wire n_4661;
wire i4_dout_606;
wire n_2216;
wire n_2206;
wire i3_dout_594;
wire n_9861;
wire n_1282;
wire n_1281;
wire n_9464;
wire n_8476;
wire n_8477;
wire n_8480;
wire n_8478;
wire u11_mem_b0_b_157;
wire n_10416;
wire n_8481;
wire n_9574;
wire oc4_int_set_716;
wire n_9575;
wire n_9450;
wire n_3341;
wire n_5683;
wire n_6163;
wire n_3278;
wire n_3000;
wire n_1323;
wire n_7933;
wire n_11462;
wire n_2237;
wire n_2387;
wire n_4568;
wire n_5463;
wire n_6137;
wire n_4569;
wire n_6136;
wire n_4632;
wire n_5454;
wire n_5791;
wire n_5278;
wire n_3982;
wire n_6132;
wire n_4603;
wire u9_mem_b1_b_131;
wire n_10309;
wire n_11097;
wire n_11100;
wire n_5676;
wire n_11099;
wire n_11098;
wire n_5670;
wire out_slt_160;
wire n_5662;
wire u10_mem_b0_b_171;
wire n_5235;
wire u11_mem_b0_b_170;
wire n_5660;
wire n_5236;
wire n_5657;
wire n_5658;
wire n_5233;
wire n_5653;
wire n_5246;
wire n_5472;
wire u10_mem_b0_b_170;
wire n_5651;
wire u11_mem_b0_b_174;
wire n_4272;
wire n_7277;
wire n_3118;
wire n_3116;
wire n_480;
wire u16_u5_dma_req_r1;
wire n_9857;
wire u10_din_tmp_53;
wire n_10095;
wire n_1012;
wire n_10329;
wire n_10404;
wire n_10405;
wire n_10085;
wire n_9990;
wire n_10094;
wire n_641;
wire n_2856;
wire in_valid_s_2;
wire n_4222;
wire n_4177;
wire n_5455;
wire n_1522;
wire n_4116;
wire n_5365;
wire n_3506;
wire n_4555;
wire n_9538;
wire n_9536;
wire n_9543;
wire o3_empty;
wire n_736;
wire n_9541;
wire n_781;
wire n_1148;
wire u11_mem_b3_b_66;
wire n_9459;
wire n_1886;
wire n_864;
wire n_7381;
wire n_7380;
wire n_8677;
wire n_1450;
wire n_7367;
wire n_4802;
wire u3_mem_b2_b_40;
wire u8_mem_b2_b_58;
wire n_1454;
wire n_7382;
wire n_7562;
wire n_10078;
wire n_12039;
wire n_4108;
wire n_2233;
wire n_2868;
wire n_2431;
wire n_3235;
wire n_1869;
wire n_2429;
wire u3_mem_b3_b_128;
wire n_10154;
wire n_1489;
wire n_8491;
wire n_10254;
wire oc2_int_set_712;
wire n_9576;
wire n_752;
wire n_683;
wire n_7276;
wire n_6324;
wire n_7135;
wire i3_dout_579;
wire n_7134;
wire i3_dout_583;
wire n_7137;
wire n_9757;
wire n_7150;
wire i3_empty;
wire n_6369;
wire n_6368;
wire u10_mem_b3_b_65;
wire n_9518;
wire n_9364;
wire n_8978;
wire n_8060;
wire n_12623;
wire u6_mem_b2_b_42;
wire u6_mem_b3_b_135;
wire u3_mem_b3_b_129;
wire n_1808;
wire u3_mem_b3_b_144;
wire u10_mem_b1_b_129;
wire n_2175;
wire n_2807;
wire n_2178;
wire n_2180;
wire n_2808;
wire n_8062;
wire n_1800;
wire u10_mem_b0_b_153;
wire n_8063;
wire n_3283;
wire n_6691;
wire n_7469;
wire n_10676;
wire n_2552;
wire n_5370;
wire n_5368;
wire n_5367;
wire n_8058;
wire u9_mem_b2_b_116;
wire n_5375;
wire n_5373;
wire n_10207;
wire n_7312;
wire n_7309;
wire n_12000;
wire n_12359;
wire n_12010;
wire n_7046;
wire n_6738;
wire n_7470;
wire n_11175;
wire u6_mem_b1_b_85;
wire n_2759;
wire n_1427;
wire n_1513;
wire n_4251;
wire n_1514;
wire u3_mem_b3_b;
wire n_1515;
wire u3_mem_b0_b_99;
wire n_10249;
wire n_9153;
wire n_8137;
wire n_10888;
wire n_6746;
wire n_612;
wire n_6747;
wire n_580;
wire n_5440;
wire n_6333;
wire n_12055;
wire n_12689;
wire n_9967;
wire n_1500;
wire n_1778;
wire n_7037;
wire n_12848;
wire n_9557;
wire n_12846;
wire n_7225;
wire n_6290;
wire n_7196;
wire n_7104;
wire n_5725;
wire n_6253;
wire n_6288;
wire n_7201;
wire n_6073;
wire n_7292;
wire n_5913;
wire n_5911;
wire n_6287;
wire n_9335;
wire n_7103;
wire n_5729;
wire n_6249;
wire n_7194;
wire n_5724;
wire n_5921;
wire n_8817;
wire n_8134;
wire u10_mem_b3_b_66;
wire n_215;
wire u10_mem_b1_b_146;
wire u11_mem_b0_b_150;
wire n_528;
wire u11_mem_b2_b_112;
wire n_12333;
wire n_12331;
wire n_8928;
wire n_2600;
wire n_4131;
wire n_3194;
wire n_4133;
wire n_4134;
wire n_3454;
wire n_3452;
wire n_6308;
wire n_4395;
wire n_6499;
wire n_6493;
wire n_6492;
wire n_10556;
wire n_5989;
wire n_10555;
wire n_6501;
wire n_10558;
wire n_6504;
wire n_5991;
wire n_6512;
wire n_10559;
wire n_6508;
wire n_3291;
wire n_1548;
wire n_6546;
wire n_8140;
wire n_8695;
wire u8_mem_b0_b_117;
wire n_3651;
wire u7_wp_b0_b;
wire n_10438;
wire u3_mem_b3_b_124;
wire n_9069;
wire n_8139;
wire n_9388;
wire n_8725;
wire n_3625;
wire n_3626;
wire n_9391;
wire n_3623;
wire n_3619;
wire n_8728;
wire u7_mem_b0_b_95;
wire n_3620;
wire n_4017;
wire n_1757;
wire n_1623;
wire n_4810;
wire n_2528;
wire n_1235;
wire n_4018;
wire n_1625;
wire n_10415;
wire n_8289;
wire n_5085;
wire n_7965;
wire n_8999;
wire n_1278;
wire n_9005;
wire n_9004;
wire n_9036;
wire n_9008;
wire n_9001;
wire n_4481;
wire n_4506;
wire n_4516;
wire n_3295;
wire n_5626;
wire n_794;
wire n_8443;
wire n_5625;
wire n_4394;
wire n_9782;
wire out_slt_103;
wire n_10951;
wire n_5492;
wire n_2326;
wire n_9975;
wire n_10674;
wire n_5293;
wire n_9519;
wire n_10354;
wire n_10353;
wire n_5490;
wire n_12018;
wire n_7175;
wire n_11676;
wire n_7199;
wire n_8175;
wire n_8673;
wire n_7440;
wire n_7384;
wire n_7385;
wire n_9456;
wire n_8177;
wire n_8674;
wire n_8181;
wire n_8675;
wire n_9458;
wire n_8178;
wire n_8676;
wire u11_mem_b0_b_166;
wire n_1263;
wire n_3784;
wire u4_mem_b0_b_108;
wire n_10633;
wire n_6227;
wire n_6225;
wire n_1001;
wire n_441;
wire n_2645;
wire n_2646;
wire n_1256;
wire n_496;
wire i6_dout_655;
wire n_4008;
wire n_457;
wire u7_wp_b2_b;
wire n_11955;
wire n_11979;
wire n_11975;
wire n_11991;
wire n_10636;
wire n_10634;
wire n_6784;
wire n_5845;
wire n_11973;
wire n_12820;
wire n_11709;
wire n_11710;
wire n_2413;
wire n_2398;
wire n_6248;
wire n_11660;
wire n_2355;
wire n_3529;
wire n_5701;
wire n_4992;
wire n_3133;
wire n_4993;
wire n_5797;
wire n_5384;
wire n_1779;
wire n_6305;
wire n_12047;
wire n_6307;
wire n_6146;
wire n_8407;
wire n_6151;
wire n_6150;
wire n_6822;
wire n_4737;
wire n_4997;
wire n_11452;
wire n_4998;
wire n_2739;
wire n_2547;
wire n_4060;
wire n_2092;
wire n_4203;
wire n_3827;
wire n_3828;
wire n_3832;
wire n_3837;
wire n_3834;
wire n_2749;
wire n_5113;
wire oc1_int_set_710;
wire n_9577;
wire n_2030;
wire n_11087;
wire n_1397;
wire n_1396;
wire n_3136;
wire n_10104;
wire u11_din_tmp_43;
wire n_10106;
wire n_4526;
wire u3_mem_b2_b_29;
wire n_1963;
wire u11_din_tmp_49;
wire u11_din_tmp_48;
wire n_4566;
wire u11_din_tmp_46;
wire n_4567;
wire u11_din_tmp_45;
wire n_8498;
wire n_8504;
wire n_8506;
wire n_8508;
wire n_8509;
wire n_8510;
wire n_6949;
wire u9_mem_b1_b_119;
wire u9_mem_b3_b_83;
wire u10_mem_b3_b_63;
wire n_4055;
wire u9_mem_b3_b_67;
wire n_11906;
wire n_6659;
wire n_6658;
wire n_6024;
wire n_5993;
wire n_6953;
wire n_6655;
wire n_6955;
wire n_6954;
wire n_6950;
wire n_6948;
wire n_6947;
wire n_2805;
wire n_2836;
wire n_3292;
wire n_8402;
wire n_8681;
wire u11_mem_b3_b_68;
wire n_10459;
wire n_6754;
wire n_7288;
wire u14_u0_full_empty_r;
wire n_9544;
wire u3_mem_b2_b_48;
wire u8_mem_b2_b;
wire n_7576;
wire n_11518;
wire n_11006;
wire n_11516;
wire n_11004;
wire n_7298;
wire n_6743;
wire u8_mem_b1_b_80;
wire n_8924;
wire n_4801;
wire n_2594;
wire n_6720;
wire n_7439;
wire n_11707;
wire n_4246;
wire n_2287;
wire n_11697;
wire n_4164;
wire n_2452;
wire u10_mem_b3_b_87;
wire n_11700;
wire n_7845;
wire u5_mem_b3_b_125;
wire n_7846;
wire u5_mem_b3_b_124;
wire n_7843;
wire n_7844;
wire n_7841;
wire n_7842;
wire n_7839;
wire u8_mem_b1_b_75;
wire n_7840;
wire n_8224;
wire n_9726;
wire n_3761;
wire n_8783;
wire n_5431;
wire n_12687;
wire n_12534;
wire n_8231;
wire u7_rp_b2_b;
wire n_9373;
wire n_11066;
wire n_8418;
wire n_8419;
wire n_7833;
wire n_8415;
wire n_4296;
wire n_7723;
wire n_8416;
wire n_7836;
wire n_8077;
wire n_4325;
wire n_8136;
wire n_8412;
wire n_8129;
wire n_4277;
wire n_8126;
wire i4_dout_614;
wire n_12521;
wire n_5378;
wire n_7702;
wire n_4635;
wire n_4792;
wire n_4636;
wire n_7701;
wire n_4595;
wire n_3555;
wire n_3914;
wire n_7704;
wire n_4389;
wire n_5058;
wire n_11988;
wire n_7230;
wire n_7079;
wire n_7203;
wire n_7081;
wire n_7227;
wire n_7306;
wire n_7271;
wire n_7095;
wire n_10504;
wire n_8213;
wire n_7285;
wire n_2595;
wire n_9580;
wire u3_mem_b1_b_80;
wire n_7695;
wire n_9131;
wire n_8475;
wire n_8173;
wire ic0_cfg_1025;
wire n_4490;
wire n_8070;
wire n_10947;
wire n_10829;
wire n_5158;
wire n_11635;
wire n_11636;
wire n_6459;
wire n_6373;
wire n_4530;
wire n_8168;
wire n_6113;
wire n_6114;
wire n_5888;
wire n_5931;
wire n_8950;
wire n_10798;
wire n_9969;
wire n_2360;
wire n_540;
wire n_10343;
wire n_9970;
wire n_10906;
wire n_7520;
wire n_565;
wire n_7434;
wire n_10799;
wire out_slt_141;
wire n_11106;
wire n_6061;
wire n_10989;
wire n_10991;
wire n_2584;
wire n_5273;
wire n_2585;
wire n_7208;
wire n_11092;
wire n_11953;
wire n_11969;
wire n_11089;
wire u9_din_tmp_51;
wire n_9788;
wire i4_dout_623;
wire n_4815;
wire n_631;
wire n_5258;
wire u13_intm_r_b8_b;
wire crac_din_699;
wire n_9434;
wire n_9125;
wire u11_mem_b2_b_96;
wire n_10476;
wire n_12377;
wire dma_req_o_b7_b;
wire n_2446;
wire n_5667;
wire n_5812;
wire n_5814;
wire n_1545;
wire n_5698;
wire n_6187;
wire n_6982;
wire n_7062;
wire n_5532;
wire n_5808;
wire n_6183;
wire n_8708;
wire n_9380;
wire n_3593;
wire n_3600;
wire n_3824;
wire n_8714;
wire n_9382;
wire u3_mem_b0_b_91;
wire n_3598;
wire n_3825;
wire n_8713;
wire n_8711;
wire n_1942;
wire n_2656;
wire n_1487;
wire n_2981;
wire n_2986;
wire n_1052;
wire n_3329;
wire n_11654;
wire n_4136;
wire n_4887;
wire n_4874;
wire n_8976;
wire n_8977;
wire n_8974;
wire u5_mem_b2_b_56;
wire n_3487;
wire oc0_cfg_964;
wire n_8555;
wire u10_mem_b3_b_80;
wire n_1723;
wire n_2655;
wire n_5129;
wire n_4497;
wire n_6613;
wire n_8522;
wire n_1716;
wire n_1715;
wire n_9926;
wire n_9927;
wire n_9928;
wire n_9929;
wire n_5870;
wire n_9922;
wire n_12836;
wire n_9925;
wire n_5866;
wire n_5864;
wire n_1807;
wire n_2696;
wire n_1938;
wire n_1939;
wire n_554;
wire u14_u5_full_empty_r;
wire n_6216;
wire n_1967;
wire n_4521;
wire n_5696;
wire n_6202;
wire n_4199;
wire n_3378;
wire n_2971;
wire n_1354;
wire n_5697;
wire n_4190;
wire n_3848;
wire n_1529;
wire n_2319;
wire n_6292;
wire n_6296;
wire n_6295;
wire n_6293;
wire n_5914;
wire n_1666;
wire n_10935;
wire n_11948;
wire n_11949;
wire n_12009;
wire n_11989;
wire n_10944;
wire n_12011;
wire n_11674;
wire n_11675;
wire n_11677;
wire n_10941;
wire n_12001;
wire n_11984;
wire n_11985;
wire n_10937;
wire n_12019;
wire u6_mem_b0_b_115;
wire n_8766;
wire u4_mem_b1_b_68;
wire n_8303;
wire n_5220;
wire n_3036;
wire n_12851;
wire n_2926;
wire n_9041;
wire n_5222;
wire n_4609;
wire n_2607;
wire n_2411;
wire n_12849;
wire n_4112;
wire n_3490;
wire n_10915;
wire oc3_int_set_713;
wire n_9784;
wire n_9785;
wire n_9786;
wire n_9868;
wire u10_din_tmp_46;
wire n_9778;
wire n_288;
wire n_10373;
wire n_129;
wire n_10382;
wire n_10383;
wire n_3213;
wire n_4551;
wire n_1915;
wire n_9233;
wire n_3866;
wire n_3411;
wire n_3082;
wire n_5169;
wire n_3074;
wire n_3066;
wire n_6506;
wire n_6067;
wire n_8485;
wire n_7458;
wire n_594;
wire u4_mem_b3_b;
wire n_8265;
wire n_2223;
wire n_2840;
wire n_11449;
wire n_1565;
wire n_9223;
wire n_2224;
wire n_2386;
wire n_1838;
wire n_2841;
wire n_12164;
wire n_8752;
wire n_9424;
wire n_9198;
wire n_7603;
wire n_7604;
wire n_10927;
wire n_5621;
wire n_4092;
wire n_3905;
wire n_9478;
wire n_8667;
wire n_7541;
wire n_8665;
wire n_9145;
wire n_11741;
wire n_12033;
wire n_3251;
wire n_3253;
wire n_3254;
wire n_11713;
wire n_2482;
wire n_11751;
wire n_5556;
wire n_6805;
wire n_11670;
wire n_11671;
wire n_4250;
wire n_6077;
wire n_1586;
wire n_1587;
wire n_4006;
wire n_1579;
wire n_9185;
wire ic1_int_set;
wire n_9485;
wire n_5003;
wire u6_mem_b1_b_80;
wire n_12355;
wire n_12358;
wire n_11842;
wire n_11844;
wire n_12125;
wire n_9108;
wire n_8373;
wire n_11015;
wire n_8088;
wire n_8107;
wire n_4324;
wire n_4293;
wire n_8397;
wire n_4480;
wire n_11178;
wire n_4896;
wire n_4895;
wire n_4894;
wire n_2715;
wire n_4900;
wire u7_mem_b1_b_76;
wire n_2706;
wire n_4899;
wire n_3103;
wire n_4897;
wire n_4891;
wire n_1430;
wire n_11738;
wire u6_mem_b3_b_141;
wire n_3177;
wire n_5050;
wire n_2802;
wire u5_mem_b1_b_69;
wire n_2760;
wire n_2717;
wire n_5045;
wire n_5044;
wire u6_mem_b3_b_139;
wire n_4383;
wire n_2051;
wire u5_mem_b1_b_72;
wire n_2725;
wire n_2785;
wire n_2535;
wire n_6610;
wire n_2537;
wire n_1672;
wire n_2536;
wire n_1671;
wire n_1215;
wire n_11623;
wire n_7118;
wire n_7211;
wire n_7059;
wire n_7210;
wire n_12062;
wire n_7215;
wire n_11627;
wire n_7119;
wire n_11994;
wire n_11901;
wire n_7213;
wire n_7060;
wire n_3956;
wire n_12843;
wire n_9960;
wire n_12809;
wire n_3668;
wire u9_mem_b2_b_103;
wire n_10280;
wire n_8823;
wire n_9052;
wire n_4433;
wire n_2052;
wire n_8301;
wire n_8017;
wire n_2047;
wire i6_dout_631;
wire n_7815;
wire n_8298;
wire n_8015;
wire n_7817;
wire n_8297;
wire n_4438;
wire n_7812;
wire n_8204;
wire n_7813;
wire n_6261;
wire n_6260;
wire n_10101;
wire n_6860;
wire n_7811;
wire u10_mem_b3_b_74;
wire n_10699;
wire n_5967;
wire n_8291;
wire n_4431;
wire n_3958;
wire n_1156;
wire n_5226;
wire n_6045;
wire n_609;
wire n_6759;
wire n_750;
wire n_541;
wire n_6671;
wire n_733;
wire n_6064;
wire n_666;
wire n_6007;
wire u10_mem_b0_b_166;
wire u11_mem_b2_b_114;
wire n_5141;
wire n_2774;
wire u10_mem_b2_b_113;
wire n_10760;
wire n_9024;
wire crac_din_695;
wire n_1034;
wire n_1524;
wire n_8184;
wire n_1229;
wire n_3521;
wire n_5881;
wire n_9806;
wire n_10919;
wire n_9807;
wire n_9808;
wire n_9810;
wire n_9811;
wire n_9812;
wire n_10926;
wire n_9813;
wire n_9815;
wire n_3132;
wire n_4623;
wire n_10441;
wire n_9804;
wire n_12835;
wire n_9376;
wire n_3746;
wire n_10130;
wire n_8692;
wire u8_mem_b0_b_121;
wire n_3822;
wire n_3748;
wire n_1732;
wire n_9371;
wire n_10812;
wire n_4524;
wire n_1703;
wire n_10466;
wire n_3523;
wire n_1252;
wire n_1251;
wire n_12584;
wire n_4957;
wire n_4931;
wire n_8955;
wire n_4909;
wire n_8954;
wire n_8958;
wire n_8956;
wire n_8960;
wire n_4862;
wire n_7634;
wire n_8959;
wire n_4959;
wire u11_mem_b1_b_119;
wire n_4618;
wire u9_din_tmp_44;
wire n_3525;
wire n_1496;
wire n_9351;
wire n_2104;
wire n_5120;
wire n_2947;
wire n_4656;
wire n_3621;
wire n_5688;
wire n_4484;
wire u3_mem_b2_b_45;
wire n_3412;
wire n_2044;
wire n_2042;
wire n_10764;
wire u14_u4_full_empty_r;
wire n_8896;
wire u10_mem_b0_b_167;
wire n_12666;
wire n_1241;
wire n_12663;
wire n_6289;
wire n_5762;
wire n_12672;
wire n_12668;
wire n_4535;
wire n_2186;
wire n_3887;
wire n_1283;
wire n_2217;
wire n_2105;
wire n_1953;
wire n_1951;
wire n_1950;
wire n_1949;
wire n_9054;
wire n_1328;
wire n_4171;
wire n_1561;
wire n_3084;
wire n_4598;
wire n_3069;
wire u11_mem_b1_b_127;
wire n_11035;
wire u11_mem_b2_b_109;
wire n_10872;
wire u11_mem_b1_b_136;
wire n_10897;
wire n_9278;
wire n_2159;
wire n_10707;
wire n_8830;
wire n_1674;
wire n_4483;
wire n_9073;
wire n_7728;
wire n_9074;
wire n_7729;
wire n_6325;
wire n_6777;
wire n_5062;
wire n_4919;
wire n_7734;
wire n_8558;
wire n_7733;
wire n_9075;
wire n_7730;
wire n_9076;
wire n_7731;
wire n_10418;
wire n_5469;
wire n_6343;
wire n_10124;
wire n_6340;
wire n_4641;
wire n_5230;
wire u10_mem_b0_b_177;
wire n_4653;
wire n_5649;
wire n_5232;
wire n_5650;
wire n_5237;
wire u10_mem_b0_b_173;
wire n_5231;
wire n_3862;
wire u9_din_tmp_45;
wire n_9775;
wire n_5644;
wire n_5234;
wire n_3875;
wire i4_dout_605;
wire n_8486;
wire n_3915;
wire n_2401;
wire n_2317;
wire n_3128;
wire n_5908;
wire n_11042;
wire n_8900;
wire u3_mem_b3_b_122;
wire u9_mem_b2_b_102;
wire u10_mem_b1_b_149;
wire n_10665;
wire n_5310;
wire n_524;
wire n_7620;
wire n_7617;
wire u3_mem_b3_b_151;
wire n_8218;
wire n_7142;
wire n_6712;
wire n_6050;
wire n_4842;
wire n_4676;
wire n_1645;
wire n_1642;
wire u11_mem_b0_b_156;
wire n_11802;
wire n_2201;
wire n_692;
wire n_2014;
wire u7_mem_b3_b_147;
wire n_2909;
wire u10_mem_b1_b_140;
wire n_5799;
wire n_5798;
wire n_8467;
wire n_6068;
wire n_7465;
wire n_10430;
wire n_8232;
wire n_6687;
wire n_7466;
wire n_8042;
wire u4_mem_b1_b_78;
wire n_5122;
wire n_8172;
wire n_4492;
wire n_8470;
wire n_4493;
wire n_8072;
wire n_2322;
wire n_863;
wire u8_mem_b2_b_55;
wire n_1871;
wire n_2902;
wire n_3364;
wire n_2029;
wire n_4323;
wire n_1974;
wire n_4911;
wire n_3258;
wire n_4429;
wire n_4386;
wire n_8792;
wire n_3656;
wire n_2212;
wire n_5090;
wire n_5089;
wire n_5092;
wire n_5091;
wire n_2941;
wire n_5087;
wire n_3293;
wire n_5086;
wire u4_mem_b3_b_145;
wire n_5088;
wire u4_mem_b3_b_143;
wire u10_mem_b0_b_160;
wire n_10135;
wire n_6251;
wire n_9638;
wire u2_bit_clk_r1;
wire i6_dout_653;
wire n_10735;
wire u9_mem_b0_b_150;
wire n_3505;
wire n_2399;
wire n_8943;
wire n_1518;
wire n_6255;
wire n_5787;
wire n_5270;
wire n_6429;
wire n_5970;
wire n_5969;
wire n_6425;
wire n_6427;
wire n_6420;
wire n_6422;
wire n_5785;
wire n_5266;
wire n_3974;
wire n_5265;
wire n_5213;
wire n_2291;
wire n_9297;
wire n_3971;
wire n_3114;
wire n_2241;
wire n_1464;
wire n_11051;
wire u11_mem_b2_b_106;
wire n_2473;
wire n_9098;
wire n_9598;
wire n_3121;
wire n_12856;
wire n_2565;
wire n_3290;
wire n_7147;
wire n_6713;
wire n_11724;
wire n_11047;
wire n_12690;
wire n_11045;
wire n_11039;
wire n_4114;
wire n_3553;
wire n_8221;
wire n_4467;
wire n_1961;
wire n_8248;
wire n_8227;
wire n_9363;
wire n_9362;
wire n_3574;
wire n_3654;
wire n_8680;
wire n_3751;
wire n_4150;
wire ic1_cfg;
wire n_2000;
wire i3_dout_593;
wire n_2489;
wire n_2962;
wire n_2961;
wire n_4126;
wire n_5619;
wire n_10301;
wire u9_mem_b3_b_60;
wire n_1651;
wire n_1648;
wire n_1162;
wire n_10867;
wire n_5311;
wire n_10868;
wire n_5322;
wire n_11109;
wire n_4244;
wire n_5316;
wire u11_mem_b2_b_97;
wire n_2022;
wire n_3086;
wire u6_mem_b0_b_114;
wire n_10625;
wire n_11104;
wire n_10953;
wire n_7530;
wire n_10622;
wire n_2669;
wire n_2668;
wire n_2665;
wire n_2667;
wire n_9151;
wire n_12683;
wire n_12686;
wire n_12682;
wire n_2663;
wire n_12685;
wire n_12116;
wire n_12684;
wire u5_mem_b0_b;
wire n_2880;
wire n_1884;
wire n_1993;
wire u9_mem_b1_b_125;
wire n_3370;
wire u8_mem_b2_b_36;
wire n_2183;
wire n_2160;
wire n_2174;
wire n_2803;
wire n_2013;
wire n_2015;
wire n_2740;
wire n_5004;
wire n_2797;
wire n_3770;
wire n_12037;
wire n_2082;
wire n_1136;
wire n_410;
wire n_11578;
wire n_5561;
wire n_5882;
wire n_37;
wire n_639;
wire n_9997;
wire n_9998;
wire n_10436;
wire n_10437;
wire n_10439;
wire n_1610;
wire n_1242;
wire n_10432;
wire n_10435;
wire n_2557;
wire n_1854;
wire n_9176;
wire n_6166;
wire n_10705;
wire n_10704;
wire n_10018;
wire n_5295;
wire n_10026;
wire n_10713;
wire n_10022;
wire n_10706;
wire n_5303;
wire n_10020;
wire n_10025;
wire n_10023;
wire u11_mem_b0_b_160;
wire u11_mem_b2_b_105;
wire n_1748;
wire u9_mem_b1_b_137;
wire n_7346;
wire n_7345;
wire n_7344;
wire n_7351;
wire n_7350;
wire n_7471;
wire n_7354;
wire i4_dout_596;
wire n_7347;
wire i4_dout_601;
wire n_7463;
wire i4_dout_602;
wire n_5865;
wire n_3193;
wire n_11440;
wire n_2438;
wire n_4814;
wire u10_mem_b0_b_152;
wire n_1891;
wire n_12810;
wire n_2560;
wire n_1337;
wire n_3288;
wire n_11655;
wire n_9546;
wire u6_mem_b3_b_126;
wire n_4638;
wire n_8447;
wire n_8448;
wire n_8450;
wire n_3843;
wire n_7985;
wire n_8442;
wire n_3874;
wire n_8152;
wire n_8437;
wire n_3880;
wire u4_mem_b3_b_137;
wire u9_mem_b1_b_120;
wire n_10300;
wire n_9174;
wire n_4039;
wire n_9426;
wire n_3285;
wire n_1986;
wire n_5094;
wire n_4925;
wire n_2946;
wire n_5098;
wire n_3305;
wire u4_mem_b3_b_135;
wire n_3844;
wire u10_mem_b3_b_59;
wire n_10566;
wire n_4922;
wire n_5097;
wire n_3434;
wire n_8049;
wire u10_mem_b1_b_128;
wire n_8487;
wire n_8435;
wire n_3881;
wire n_8149;
wire u9_mem_b1_b_134;
wire n_10305;
wire n_7165;
wire n_7712;
wire n_9749;
wire n_1972;
wire n_8426;
wire n_2157;
wire u10_mem_b3_b_64;
wire n_8815;
wire n_2152;
wire n_2766;
wire n_3279;
wire n_3280;
wire u7_mem_b3_b_143;
wire n_3535;
wire n_8932;
wire n_605;
wire n_2370;
wire n_6461;
wire n_6464;
wire n_6467;
wire n_6455;
wire n_6243;
wire n_5875;
wire n_6451;
wire n_3076;
wire n_3764;
wire u4_mem_b0_b_117;
wire n_3763;
wire u5_mem_b2_b_47;
wire n_12050;
wire n_4224;
wire n_3437;
wire n_1794;
wire n_549;
wire n_543;
wire n_12049;
wire n_12056;
wire n_3557;
wire n_12053;
wire n_3424;
wire n_8523;
wire n_8525;
wire n_8530;
wire n_8532;
wire n_2457;
wire n_5595;
wire n_4601;
wire n_2923;
wire n_340;
wire u9_mem_b1_b_126;
wire n_1793;
wire n_557;
wire n_574;
wire n_12077;
wire n_10302;
wire n_6885;
wire n_1243;
wire n_10984;
wire n_1885;
wire n_11064;
wire n_11065;
wire n_10619;
wire n_11068;
wire n_9130;
wire u9_mem_b2_b_92;
wire u5_mem_b2_b_44;
wire n_2879;
wire n_2883;
wire u11_mem_b3_b_67;
wire n_3780;
wire n_9211;
wire n_743;
wire u11_mem_b3_b_64;
wire n_10655;
wire n_3779;
wire u4_mem_b0_b_110;
wire n_12804;
wire n_257;
wire n_1105;
wire n_1185;
wire n_2357;
wire n_2478;
wire n_3776;
wire n_974;
wire n_197;
wire n_4034;
wire n_3773;
wire n_12735;
wire n_1975;
wire n_4503;
wire n_3151;
wire n_2199;
wire n_3425;
wire n_5134;
wire n_2905;
wire n_10472;
wire n_10809;
wire n_10830;
wire n_10409;
wire n_10966;
wire oc1_int_set;
wire n_10832;
wire n_610;
wire n_11009;
wire n_10808;
wire n_10407;
wire n_1037;
wire n_1746;
wire n_1747;
wire n_4617;
wire n_3416;
wire n_4605;
wire n_7770;
wire n_4545;
wire n_7773;
wire n_9128;
wire n_4543;
wire n_4358;
wire n_4547;
wire n_7772;
wire n_9129;
wire n_5156;
wire n_4851;
wire n_3407;
wire u3_mem_b1_b_87;
wire n_2769;
wire n_7377;
wire n_1022;
wire n_3981;
wire n_7157;
wire n_7294;
wire n_7032;
wire n_10458;
wire n_10083;
wire n_5079;
wire n_2588;
wire n_2575;
wire u11_mem_b0_b_159;
wire n_8925;
wire n_9992;
wire n_10392;
wire n_312;
wire n_9497;
wire n_9486;
wire n_9559;
wire n_9548;
wire n_9498;
wire n_9488;
wire u9_mem_b2_b_89;
wire n_9558;
wire n_3150;
wire i4_empty;
wire n_8639;
wire u10_mem_b2_b_106;
wire n_5581;
wire n_5583;
wire n_5743;
wire n_5161;
wire n_5740;
wire n_5738;
wire u10_mem_b0_b;
wire u11_mem_b2_b_115;
wire n_10052;
wire n_206;
wire n_10053;
wire n_12157;
wire n_6200;
wire n_3027;
wire n_12841;
wire n_12855;
wire n_12798;
wire n_5562;
wire n_1506;
wire n_9155;
wire n_5899;
wire n_8827;
wire n_9439;
wire u4_mem_b0_b_109;
wire n_3783;
wire n_8822;
wire n_8944;
wire i4_dout_615;
wire n_9229;
wire n_9102;
wire n_7998;
wire n_7999;
wire n_8000;
wire n_8001;
wire n_7444;
wire u5_mem_b3_b_123;
wire n_9209;
wire u8_mem_b3_b_145;
wire n_8852;
wire n_4061;
wire u5_mem_b2_b_33;
wire n_4923;
wire n_3410;
wire n_8599;
wire n_8796;
wire n_4327;
wire n_1806;
wire n_9045;
wire n_10840;
wire n_4338;
wire n_2080;
wire n_4932;
wire n_4934;
wire n_2838;
wire n_1273;
wire n_1996;
wire n_8909;
wire n_9067;
wire n_4867;
wire n_7589;
wire n_8127;
wire n_7721;
wire n_9066;
wire n_7722;
wire n_5308;
wire n_5318;
wire n_8122;
wire n_5314;
wire n_5323;
wire u11_mem_b1_b_139;
wire n_8282;
wire i6_dout_630;
wire n_5869;
wire n_5871;
wire n_8283;
wire n_5873;
wire n_2609;
wire n_1776;
wire u4_mem_b2_b_59;
wire n_8273;
wire n_7948;
wire n_8121;
wire u5_mem_b2_b_55;
wire n_9252;
wire u4_mem_b0_b_119;
wire n_8818;
wire n_7799;
wire n_7798;
wire n_3617;
wire n_12058;
wire n_3910;
wire n_4573;
wire n_2462;
wire n_3054;
wire n_5199;
wire n_4159;
wire n_3051;
wire n_8566;
wire n_8563;
wire oc1_cfg_980;
wire n_8562;
wire n_1076;
wire n_10856;
wire n_3615;
wire n_6889;
wire n_6888;
wire n_10281;
wire n_6874;
wire n_10276;
wire n_10275;
wire n_2236;
wire n_2479;
wire n_2908;
wire n_3940;
wire n_11533;
wire n_127;
wire n_453;
wire oc1_cfg;
wire n_1132;
wire n_8410;
wire n_2327;
wire u15_valid_r;
wire n_3302;
wire n_12156;
wire n_6741;
wire n_597;
wire u9_mem_b3_b_87;
wire n_10700;
wire n_9720;
wire n_447;
wire n_9705;
wire n_5585;
wire n_4733;
wire n_5680;
wire n_1200;
wire n_8901;
wire n_2483;
wire n_553;
wire n_12751;
wire n_656;
wire n_8765;
wire u3_mem_b1_b_73;
wire n_8767;
wire n_9407;
wire n_3614;
wire n_8760;
wire u11_mem_b3_b_79;
wire n_10853;
wire u10_mem_b3_b_81;
wire n_4341;
wire n_7286;
wire n_10757;
wire n_10833;
wire n_11014;
wire n_11012;
wire n_10831;
wire n_4631;
wire n_3554;
wire n_3939;
wire n_709;
wire n_10864;
wire n_4630;
wire n_2461;
wire n_2640;
wire n_9101;
wire n_9100;
wire n_7750;
wire n_9060;
wire n_9106;
wire n_4924;
wire n_7754;
wire n_7748;
wire n_7749;
wire n_10740;
wire n_3970;
wire n_6997;
wire n_7115;
wire n_5880;
wire n_3968;
wire n_3969;
wire u13_ints_r_b9_b;
wire n_3966;
wire n_8751;
wire u14_u1_full_empty_r;
wire n_9542;
wire o3_status_962;
wire n_1899;
wire n_8304;
wire n_3893;
wire ic1_int_set_722;
wire u9_mem_b3_b;
wire n_10049;
wire n_10050;
wire n_10047;
wire n_1863;
wire n_10048;
wire n_10044;
wire n_10046;
wire n_10042;
wire n_35;
wire n_10043;
wire n_9183;
wire n_416;
wire n_4762;
wire n_4760;
wire n_10766;
wire n_5416;
wire u11_mem_b0_b_168;
wire n_5415;
wire n_5414;
wire n_5412;
wire u9_mem_b0_b_163;
wire n_8310;
wire n_3060;
wire n_1326;
wire n_1542;
wire n_8236;
wire n_8849;
wire n_8067;
wire n_4856;
wire n_7563;
wire n_2280;
wire n_7869;
wire n_11924;
wire n_8018;
wire n_8229;
wire n_8019;
wire n_8020;
wire n_8022;
wire n_8023;
wire n_7946;
wire n_7445;
wire u3_mem_b1_b_79;
wire n_8812;
wire n_1707;
wire n_11034;
wire n_2279;
wire n_10098;
wire n_2332;
wire n_12063;
wire n_11628;
wire n_11995;
wire n_6185;
wire n_11618;
wire n_11620;
wire n_11624;
wire n_10224;
wire u6_wp_b0_b;
wire n_4945;
wire n_2737;
wire n_4944;
wire n_2787;
wire oc2_cfg;
wire n_4427;
wire n_1991;
wire n_5111;
wire n_2102;
wire n_2682;
wire n_1976;
wire n_2690;
wire n_5114;
wire n_6334;
wire u7_mem_b3_b_142;
wire n_10119;
wire n_5946;
wire n_2123;
wire n_8780;
wire n_3328;
wire n_2384;
wire n_3741;
wire n_8902;
wire n_2290;
wire n_3111;
wire n_11922;
wire n_11928;
wire n_3112;
wire n_1536;
wire n_5211;
wire n_3173;
wire n_3563;
wire n_8589;
wire ic2_cfg_1050;
wire n_8597;
wire n_6583;
wire n_6921;
wire n_6608;
wire n_6923;
wire n_10252;
wire n_10247;
wire n_6892;
wire u10_mem_b0_b_165;
wire n_4858;
wire u3_mem_b1_b_82;
wire n_11501;
wire n_10666;
wire n_4673;
wire n_5481;
wire n_2937;
wire u10_mem_b0_b_155;
wire n_1335;
wire n_5708;
wire i6_dout_650;
wire i4_dout_624;
wire n_10097;
wire n_3422;
wire n_3420;
wire n_9277;
wire n_9419;
wire n_8782;
wire n_9416;
wire n_3820;
wire n_968;
wire n_412;
wire n_9774;
wire n_4807;
wire n_9276;
wire n_4972;
wire n_4973;
wire n_2821;
wire n_4970;
wire n_4971;
wire n_4976;
wire n_4974;
wire n_4975;
wire n_1702;
wire n_4968;
wire n_4969;
wire n_9173;
wire u11_mem_b2_b_104;
wire n_10841;
wire n_9867;
wire n_4670;
wire n_3363;
wire n_4671;
wire n_4672;
wire n_2895;
wire n_2576;
wire u9_mem_b1_b_129;
wire n_8490;
wire n_5436;
wire n_12481;
wire n_6218;
wire n_6778;
wire u9_mem_b2_b_96;
wire n_10014;
wire n_10015;
wire u9_mem_b3_b_74;
wire n_10016;
wire n_10017;
wire n_10728;
wire i3_dout_570;
wire n_10739;
wire n_10732;
wire n_8215;
wire n_5400;
wire n_8264;
wire n_9578;
wire n_6667;
wire n_6666;
wire n_6669;
wire n_6611;
wire n_6036;
wire n_10326;
wire n_5999;
wire n_10657;
wire n_10659;
wire n_3181;
wire n_2298;
wire n_2299;
wire n_7574;
wire n_8878;
wire n_4559;
wire n_2274;
wire n_4158;
wire n_4157;
wire n_7968;
wire n_7442;
wire n_4958;
wire n_7966;
wire n_5142;
wire n_12167;
wire n_12617;
wire n_8641;
wire u14_u2_full_empty_r;
wire n_9539;
wire n_12618;
wire n_12611;
wire n_9607;
wire n_6709;
wire n_869;
wire n_7978;
wire n_7986;
wire n_7851;
wire n_1532;
wire n_3754;
wire n_3756;
wire n_3757;
wire n_4416;
wire n_2089;
wire u4_mem_b2_b_33;
wire n_3762;
wire n_2754;
wire n_2172;
wire n_7724;
wire n_2097;
wire n_5029;
wire n_5031;
wire n_5030;
wire n_2771;
wire n_10877;
wire n_3753;
wire n_604;
wire n_4712;
wire n_4715;
wire n_4709;
wire n_4707;
wire n_8635;
wire n_8633;
wire n_8638;
wire n_8637;
wire n_8630;
wire n_6580;
wire n_6587;
wire n_6015;
wire n_6012;
wire n_6009;
wire n_10232;
wire n_10230;
wire n_6593;
wire n_5861;
wire n_7100;
wire n_7101;
wire n_5717;
wire n_6240;
wire n_5858;
wire n_9338;
wire n_9433;
wire n_2873;
wire u9_mem_b3_b_58;
wire n_3007;
wire n_7372;
wire n_7374;
wire n_7153;
wire n_7152;
wire n_2407;
wire i3_dout_566;
wire n_11668;
wire n_997;
wire n_3409;
wire n_1492;
wire n_1728;
wire u9_mem_b0_b_176;
wire n_8803;
wire n_8798;
wire n_8800;
wire u5_mem_b0_b_91;
wire n_3724;
wire u8_mem_b3_b_142;
wire n_8203;
wire valid_s1;
wire n_1750;
wire n_9535;
wire n_1711;
wire n_4558;
wire n_1901;
wire n_4988;
wire n_2987;
wire n_4989;
wire n_4990;
wire n_4268;
wire n_11450;
wire n_4267;
wire n_4269;
wire n_7789;
wire n_4468;
wire n_7790;
wire n_10898;
wire n_7792;
wire n_7793;
wire n_9150;
wire n_7794;
wire n_7795;
wire u9_mem_b0_b_164;
wire n_8403;
wire n_2140;
wire u11_mem_b2_b_118;
wire n_8654;
wire n_10818;
wire n_1258;
wire n_5394;
wire n_4068;
wire n_10890;
wire n_9525;
wire n_9840;
wire n_9599;
wire n_8905;
wire n_7593;
wire n_7594;
wire n_8124;
wire n_8903;
wire n_3841;
wire n_7590;
wire n_7591;
wire n_8897;
wire n_7725;
wire n_7726;
wire n_8895;
wire n_4275;
wire n_7586;
wire n_4274;
wire n_7587;
wire u10_mem_b1_b_127;
wire n_6458;
wire n_10521;
wire n_5979;
wire n_5978;
wire n_10514;
wire n_5995;
wire n_1204;
wire u5_mem_b2_b_57;
wire n_11476;
wire u5_mem_b2_b_45;
wire i6_dout_628;
wire i6_dout_629;
wire i3_dout_592;
wire n_839;
wire n_1174;
wire n_4824;
wire n_8064;
wire n_2173;
wire n_4470;
wire n_1792;
wire n_4469;
wire n_4463;
wire n_4465;
wire n_1741;
wire n_4462;
wire n_9521;
wire suspended_o;
wire n_830;
wire n_2087;
wire n_3210;
wire n_9484;
wire n_3208;
wire n_2210;
wire n_4637;
wire n_3946;
wire n_9021;
wire n_1846;
wire n_9204;
wire n_7849;
wire n_9208;
wire n_7848;
wire n_9207;
wire n_7847;
wire n_9206;
wire n_5679;
wire n_4380;
wire n_2373;
wire n_8935;
wire n_5255;
wire n_4694;
wire n_4693;
wire n_4692;
wire n_9063;
wire n_4689;
wire n_8929;
wire n_569;
wire n_2810;
wire n_4093;
wire n_5887;
wire n_5883;
wire n_5885;
wire n_5878;
wire n_10827;
wire u10_mem_b2_b_103;
wire n_1512;
wire n_1883;
wire n_1090;
wire n_2392;
wire u11_din_tmp_44;
wire n_10102;
wire n_4817;
wire n_2393;
wire u11_mem_b0_b_165;
wire n_2221;
wire n_2839;
wire n_2215;
wire u13_ints_r_b13_b;
wire n_1865;
wire n_6604;
wire n_4217;
wire n_3394;
wire n_12833;
wire n_3760;
wire n_8813;
wire n_7868;
wire n_7867;
wire u10_mem_b3_b_76;
wire u8_mem_b3_b_129;
wire n_4994;
wire n_2939;
wire n_3234;
wire n_4362;
wire n_4363;
wire n_4360;
wire n_4361;
wire n_4357;
wire n_9827;
wire n_12374;
wire n_9257;
wire n_11499;
wire n_4608;
wire n_5528;
wire n_2382;
wire n_6188;
wire u11_mem_b3_b_82;
wire n_8305;
wire n_719;
wire n_4054;
wire n_1749;
wire n_1752;
wire n_1751;
wire n_12048;
wire n_1759;
wire n_1758;
wire n_1753;
wire n_9231;
wire n_9452;
wire n_10773;
wire n_10332;
wire n_12256;
wire n_10331;
wire n_10774;
wire n_9963;
wire n_9547;
wire n_9586;
wire n_9482;
wire n_9585;
wire n_10776;
wire n_8922;
wire n_4282;
wire u11_mem_b3_b_58;
wire n_6605;
wire n_10462;
wire n_6555;
wire n_10837;
wire n_7882;
wire n_7883;
wire n_8750;
wire n_8411;
wire n_7886;
wire n_7887;
wire n_8479;
wire n_7885;
wire n_6055;
wire n_4035;
wire n_8367;
wire n_2837;
wire n_11176;
wire n_9693;
wire n_9692;
wire n_7934;
wire n_7935;
wire n_2337;
wire n_5716;
wire n_7932;
wire n_9741;
wire n_5715;
wire n_4447;
wire n_4446;
wire n_12853;
wire n_12854;
wire n_3867;
wire n_4450;
wire n_4449;
wire n_4448;
wire n_5115;
wire n_4451;
wire n_11112;
wire n_12032;
wire oc1_int_set_709;
wire u9_mem_b2_b_97;
wire n_1511;
wire n_4207;
wire n_9834;
wire n_9686;
wire n_9533;
wire n_5299;
wire n_5305;
wire n_8821;
wire n_2943;
wire n_7269;
wire n_6998;
wire n_2633;
wire n_2813;
wire u10_mem_b0_b_157;
wire n_6974;
wire n_6969;
wire n_6971;
wire n_6975;
wire n_5567;
wire n_6082;
wire n_7052;
wire n_5572;
wire n_6967;
wire n_6968;
wire n_1030;
wire n_8468;
wire n_8187;
wire n_8285;
wire n_2453;
wire u10_mem_b3_b_68;
wire n_9281;
wire wb_ack_o;
wire n_9064;
wire n_2197;
wire n_2261;
wire n_3898;
wire n_3896;
wire n_2472;
wire n_2296;
wire n_2820;
wire n_5819;
wire n_6199;
wire u9_mem_b1_b_123;
wire n_1347;
wire n_1646;
wire n_1640;
wire n_6976;
wire n_10894;
wire n_9569;
wire n_928;
wire n_6557;
wire n_10178;
wire n_10825;
wire n_2264;
wire n_4040;
wire n_7994;
wire n_11651;
wire n_1142;
wire n_4178;
wire n_4600;
wire n_12536;
wire n_11181;
wire n_6043;
wire n_9850;
wire n_10355;
wire n_7162;
wire n_6996;
wire n_6993;
wire n_7102;
wire n_2940;
wire n_5790;
wire n_2198;
wire n_2167;
wire n_865;
wire n_6750;
wire n_1000;
wire n_8306;
wire n_8302;
wire n_4295;
wire n_1259;
wire n_1289;
wire n_12803;
wire n_3126;
wire n_2894;
wire n_11460;
wire n_4301;
wire n_7890;
wire n_7889;
wire n_7888;
wire n_9249;
wire n_5275;
wire n_4725;
wire n_3991;
wire u9_mem_b0_b_152;
wire i4_dout_612;
wire n_5391;
wire n_9299;
wire n_10156;
wire n_7910;
wire n_7909;
wire n_7912;
wire n_7911;
wire u9_mem_b1_b_128;
wire n_8489;
wire n_9339;
wire n_2906;
wire n_12372;
wire u9_mem_b1_b;
wire n_5726;
wire n_12365;
wire n_4239;
wire n_3195;
wire n_8109;
wire n_1143;
wire n_5364;
wire n_10695;
wire n_5521;
wire n_10697;
wire n_5366;
wire n_10703;
wire n_5517;
wire n_5519;
wire n_12168;
wire oc0_int_set;
wire n_5479;
wire n_5482;
wire n_5483;
wire n_5475;
wire n_5477;
wire n_10151;
wire n_5473;
wire i4_dout_611;
wire n_8330;
wire n_1231;
wire n_5860;
wire n_5776;
wire n_7268;
wire n_5775;
wire n_7270;
wire n_5757;
wire n_7319;
wire n_7273;
wire n_6125;
wire n_4342;
wire n_3376;
wire n_5392;
wire n_10675;
wire n_9451;
wire n_2907;
wire n_8167;
wire n_8048;
wire n_8342;
wire n_8052;
wire n_6973;
wire n_9280;
wire n_4379;
wire n_7698;
wire n_4376;
wire n_4375;
wire n_7699;
wire n_9042;
wire u11_mem_b2_b_94;
wire n_7703;
wire n_3342;
wire n_2858;
wire n_8186;
wire n_8185;
wire n_2998;
wire n_6095;
wire n_5539;
wire n_6097;
wire n_5456;
wire n_6099;
wire n_5457;
wire n_6761;
wire n_5699;
wire n_5756;
wire n_4154;
wire n_12496;
wire n_12495;
wire n_9304;
wire n_4806;
wire n_3013;
wire dma_req_o_b5_b;
wire n_8496;
wire out_slt6;
wire n_10952;
wire out_slt_122;
wire n_11110;
wire n_7021;
wire n_3701;
wire n_3037;
wire n_8404;
wire n_10858;
wire n_10819;
wire n_745;
wire n_1197;
wire n_8809;
wire n_9977;
wire n_9978;
wire n_10357;
wire n_10358;
wire n_5362;
wire n_9976;
wire n_5495;
wire n_10356;
wire n_5491;
wire n_5349;
wire i4_dout_595;
wire n_587;
wire n_10133;
wire n_10138;
wire n_11659;
wire n_11913;
wire n_11911;
wire n_11927;
wire u11_mem_b1_b_132;
wire n_6108;
wire n_6109;
wire n_8753;
wire n_12832;
wire n_5587;
wire n_1189;
wire n_11465;
wire n_3918;
wire n_7138;
wire n_5590;
wire n_7139;
wire n_5789;
wire n_4118;
wire n_5686;
wire n_4660;
wire n_4664;
wire n_4663;
wire n_9298;
wire n_12378;
wire out_slt8;
wire n_11107;
wire n_12480;
wire n_3098;
wire n_5459;
wire n_12478;
wire oc2_cfg_989;
wire n_7481;
wire n_9401;
wire u10_mem_b3_b_83;
wire n_9344;
wire n_700;
wire n_10863;
wire n_7447;
wire n_7449;
wire n_10954;
wire n_10950;
wire n_9987;
wire u9_mem_b3_b_63;
wire u14_n_135;
wire out_slt3;
wire n_11103;
wire u11_mem_b2_b_102;
wire n_12829;
wire n_12830;
wire n_1997;
wire n_10399;
wire n_5910;
wire n_2511;
wire n_2359;
wire n_3895;
wire n_8284;
wire n_7568;
wire n_7719;
wire n_2872;
wire n_10100;
wire oc5_cfg;
wire n_11987;
wire n_12457;
wire n_12458;
wire n_6286;
wire n_5474;
wire n_11669;
wire n_11703;
wire n_3109;
wire n_2874;
wire n_11704;
wire n_9572;
wire n_11897;
wire n_11900;
wire n_9776;
wire n_4347;
wire n_6994;
wire n_7173;
wire n_8488;
wire n_12114;
wire n_1159;
wire n_8123;
wire n_3287;
wire n_2999;
wire n_1348;
wire n_9340;
wire n_1910;
wire n_11108;
wire n_2510;
wire n_2859;
wire n_846;
// scan chain begins here
SDFFN u16_u1_dma_req_reg (.CK(clk_i), .D(n_11194), .Q(dma_req_o_b1_b), .SO(dma_req_o_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(scan_data_in));
SDFFN u16_u3_dma_req_reg (.CK(clk_i), .D(n_11193), .Q(dma_req_o_b3_b), .SO(dma_req_o_b3_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(dma_req_o_b1_b));
SDFFN u16_u0_dma_req_reg (.CK(clk_i), .D(n_11192), .Q(dma_req_o_b0_b), .SO(dma_req_o_b0_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(dma_req_o_b3_b));
SDFFN u16_u2_dma_req_reg (.CK(clk_i), .D(n_11191), .Q(dma_req_o_b2_b), .SO(dma_req_o_b2_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(dma_req_o_b0_b));
SDFFN u16_u4_dma_req_reg (.CK(clk_i), .D(n_11190), .Q(dma_req_o_b4_b), .SO(dma_req_o_b4_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(dma_req_o_b2_b));
SDFFN u16_u5_dma_req_reg (.CK(clk_i), .D(n_11189), .Q(dma_req_o_b5_b), .SO(dma_req_o_b5_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(dma_req_o_b4_b));
SDFFN u4_rp_reg_b2_b (.CK(clk_i), .D(n_11165), .Q(u4_rp_b2_b), .SO(u4_rp_b2_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(dma_req_o_b5_b));
SDFFN u5_rp_reg_b2_b (.CK(clk_i), .D(n_11164), .Q(u5_rp_b2_b), .SO(u5_rp_b2_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_rp_b2_b));
SDFFN u8_rp_reg_b2_b (.CK(clk_i), .D(n_11181), .Q(u8_rp_b2_b), .SO(u8_rp_b2_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_rp_b2_b));
SDFFN u3_rp_reg_b2_b (.CK(clk_i), .D(n_11180), .Q(u3_rp_b2_b), .SO(u3_rp_b2_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_rp_b2_b));
SDFFN u6_rp_reg_b2_b (.CK(clk_i), .D(n_11179), .Q(u6_rp_b2_b), .SO(u6_rp_b2_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_rp_b2_b));
SDFFN u7_rp_reg_b2_b (.CK(clk_i), .D(n_11178), .Q(u7_rp_b2_b), .SO(u7_rp_b2_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_rp_b2_b));
SDFFN u8_rp_reg_b3_b (.CK(clk_i), .D(n_12592), .Q(u8_rp_b3_b), .SO(u8_rp_b3_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_rp_b2_b));
SDFFN u3_rp_reg_b3_b (.CK(clk_i), .D(n_11176), .Q(u3_rp_b3_b), .SO(u3_rp_b3_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_rp_b3_b));
SDFFN u6_rp_reg_b3_b (.CK(clk_i), .D(n_11175), .Q(u6_rp_b3_b), .SO(u6_rp_b3_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_rp_b3_b));
SDFFN u7_rp_reg_b3_b (.CK(clk_i), .D(n_11174), .Q(u7_rp_b3_b), .SO(u7_rp_b3_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_rp_b3_b));
SDFFN u8_rp_reg_b1_b (.CK(clk_i), .D(n_11163), .Q(u8_rp_b1_b), .SO(u8_rp_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_rp_b3_b));
SDFFN u3_rp_reg_b1_b (.CK(clk_i), .D(n_11162), .Q(u3_rp_b1_b), .SO(u3_rp_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_rp_b1_b));
SDFFN u7_rp_reg_b1_b (.CK(clk_i), .D(n_11160), .Q(u7_rp_b1_b), .SO(u7_rp_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_rp_b1_b));
SDFFN u6_rp_reg_b1_b (.CK(clk_i), .D(n_11161), .Q(u6_rp_b1_b), .SO(u6_rp_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_rp_b1_b));
SDFFN u13_ints_r_reg_b11_b (.CK(clk_i), .D(n_11121), .Q(u13_ints_r_b11_b), .SO(u13_ints_r_b11_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_rp_b1_b));
SDFFN u13_ints_r_reg_b5_b (.CK(clk_i), .D(n_11120), .Q(u13_ints_r_b5_b), .SO(u13_ints_r_b5_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b11_b));
SDFFN u4_rp_reg_b1_b (.CK(clk_i), .D(n_11153), .Q(u4_rp_b1_b), .SO(u4_rp_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b5_b));
SDFFN u4_rp_reg_b3_b (.CK(clk_i), .D(n_11157), .Q(u4_rp_b3_b), .SO(u4_rp_b3_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_rp_b1_b));
SDFFN u5_rp_reg_b1_b (.CK(clk_i), .D(n_11152), .Q(u5_rp_b1_b), .SO(u5_rp_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_rp_b3_b));
SDFFN u5_rp_reg_b3_b (.CK(clk_i), .D(n_11155), .Q(u5_rp_b3_b), .SO(u5_rp_b3_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_rp_b1_b));
SDFFNSRN u6_dout_reg_b2_b (.CK(clk_i), .D(n_11149), .Q(out_slt_123), .SO(out_slt_123), .SE(scan_enable), .SI(u5_rp_b3_b));
SDFFNSRN u6_dout_reg_b3_b (.CK(clk_i), .D(n_11148), .Q(out_slt_124), .SO(out_slt_124), .SE(scan_enable), .SI(out_slt_123));
SDFFNSRN u7_dout_reg_b2_b (.CK(clk_i), .D(n_11146), .Q(out_slt_142), .SO(out_slt_142), .SE(scan_enable), .SI(out_slt_124));
SDFFNSRN u7_dout_reg_b3_b (.CK(clk_i), .D(n_11145), .Q(out_slt_143), .SO(out_slt_143), .SE(scan_enable), .SI(out_slt_142));
SDFFNSRN u3_dout_reg_b2_b (.CK(clk_i), .D(n_11135), .Q(out_slt_66), .SO(out_slt_66), .SE(scan_enable), .SI(out_slt_143));
SDFFNSRN u3_dout_reg_b3_b (.CK(clk_i), .D(n_11134), .Q(out_slt_67), .SO(out_slt_67), .SE(scan_enable), .SI(out_slt_66));
SDFFNSRN u8_dout_reg_b2_b (.CK(clk_i), .D(n_11130), .Q(out_slt_161), .SO(out_slt_161), .SE(scan_enable), .SI(out_slt_67));
SDFFNSRN u8_dout_reg_b3_b (.CK(clk_i), .D(n_11129), .Q(out_slt_162), .SO(out_slt_162), .SE(scan_enable), .SI(out_slt_161));
SDFFN u13_ints_r_reg_b14_b (.CK(clk_i), .D(n_11015), .Q(u13_ints_r_b14_b), .SO(u13_ints_r_b14_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(out_slt_162));
SDFFN u13_ints_r_reg_b17_b (.CK(clk_i), .D(n_11014), .Q(u13_ints_r_b17_b), .SO(u13_ints_r_b17_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b14_b));
SDFFN u13_ints_r_reg_b2_b (.CK(clk_i), .D(n_11012), .Q(u13_ints_r_b2_b), .SO(u13_ints_r_b2_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b17_b));
SDFFN u13_ints_r_reg_b8_b (.CK(clk_i), .D(n_11011), .Q(u13_ints_r_b8_b), .SO(u13_ints_r_b8_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b2_b));
SDFFNSRN u6_dout_reg_b0_b (.CK(clk_i), .D(n_11111), .Q(out_slt7), .SO(out_slt7), .SE(scan_enable), .SI(u13_ints_r_b8_b));
SDFFNSRN u6_dout_reg_b1_b (.CK(clk_i), .D(n_11110), .Q(out_slt_122), .SO(out_slt_122), .SE(scan_enable), .SI(out_slt7));
SDFFNSRN u7_dout_reg_b0_b (.CK(clk_i), .D(n_11107), .Q(out_slt8), .SO(out_slt8), .SE(scan_enable), .SI(out_slt_122));
SDFFNSRN u7_dout_reg_b1_b (.CK(clk_i), .D(n_11106), .Q(out_slt_141), .SO(out_slt_141), .SE(scan_enable), .SI(out_slt8));
SDFFNSRN u3_dout_reg_b0_b (.CK(clk_i), .D(n_11103), .Q(out_slt3), .SO(out_slt3), .SE(scan_enable), .SI(out_slt_141));
SDFFNSRN u8_dout_reg_b0_b (.CK(clk_i), .D(n_11102), .Q(out_slt9), .SO(out_slt9), .SE(scan_enable), .SI(out_slt3));
SDFFNSRN u3_dout_reg_b1_b (.CK(clk_i), .D(n_11101), .Q(out_slt_65), .SO(out_slt_65), .SE(scan_enable), .SI(out_slt9));
SDFFNSRN u8_dout_reg_b1_b (.CK(clk_i), .D(n_11098), .Q(out_slt_160), .SO(out_slt_160), .SE(scan_enable), .SI(out_slt_65));
SDFFNSRN u8_rp_reg_b0_b (.CK(clk_i), .D(n_11009), .Q(n_610), .SO(n_610), .SE(scan_enable), .SI(out_slt_160));
SDFFNSRN u3_rp_reg_b0_b (.CK(clk_i), .D(n_11008), .Q(u3_rp_b0_b), .SO(u3_rp_b0_b), .SE(scan_enable), .SI(n_610));
SDFFNSRN u6_rp_reg_b0_b (.CK(clk_i), .D(n_11113), .Q(u6_rp_b0_b), .SO(u6_rp_b0_b), .SE(scan_enable), .SI(u3_rp_b0_b));
SDFFNSRN u7_rp_reg_b0_b (.CK(clk_i), .D(n_11112), .Q(u7_rp_b0_b), .SO(u7_rp_b0_b), .SE(scan_enable), .SI(u6_rp_b0_b));
SDFFNSRN u6_dout_reg_b12_b (.CK(clk_i), .D(n_11093), .Q(out_slt_133), .SO(out_slt_133), .SE(scan_enable), .SI(u7_rp_b0_b));
SDFFNSRN u6_dout_reg_b13_b (.CK(clk_i), .D(n_11092), .Q(out_slt_134), .SO(out_slt_134), .SE(scan_enable), .SI(out_slt_133));
SDFFNSRN u6_dout_reg_b14_b (.CK(clk_i), .D(n_11091), .Q(out_slt_135), .SO(out_slt_135), .SE(scan_enable), .SI(out_slt_134));
SDFFNSRN u6_dout_reg_b15_b (.CK(clk_i), .D(n_11089), .Q(out_slt_136), .SO(out_slt_136), .SE(scan_enable), .SI(out_slt_135));
SDFFNSRN u6_dout_reg_b10_b (.CK(clk_i), .D(n_11095), .Q(out_slt_131), .SO(out_slt_131), .SE(scan_enable), .SI(out_slt_136));
SDFFNSRN u6_dout_reg_b11_b (.CK(clk_i), .D(n_11094), .Q(out_slt_132), .SO(out_slt_132), .SE(scan_enable), .SI(out_slt_131));
SDFFNSRN u6_dout_reg_b18_b (.CK(clk_i), .D(n_11084), .Q(out_slt_139), .SO(out_slt_139), .SE(scan_enable), .SI(out_slt_132));
SDFFNSRN u6_dout_reg_b19_b (.CK(clk_i), .D(n_11082), .Q(out_slt_140), .SO(out_slt_140), .SE(scan_enable), .SI(out_slt_139));
SDFFNSRN u6_dout_reg_b16_b (.CK(clk_i), .D(n_11087), .Q(out_slt_137), .SO(out_slt_137), .SE(scan_enable), .SI(out_slt_140));
SDFFNSRN u6_dout_reg_b17_b (.CK(clk_i), .D(n_11085), .Q(out_slt_138), .SO(out_slt_138), .SE(scan_enable), .SI(out_slt_137));
SDFFNSRN u6_dout_reg_b4_b (.CK(clk_i), .D(n_11081), .Q(out_slt_125), .SO(out_slt_125), .SE(scan_enable), .SI(out_slt_138));
SDFFNSRN u6_dout_reg_b5_b (.CK(clk_i), .D(n_11080), .Q(out_slt_126), .SO(out_slt_126), .SE(scan_enable), .SI(out_slt_125));
SDFFNSRN u6_dout_reg_b6_b (.CK(clk_i), .D(n_11079), .Q(out_slt_127), .SO(out_slt_127), .SE(scan_enable), .SI(out_slt_126));
SDFFNSRN u6_dout_reg_b7_b (.CK(clk_i), .D(n_11078), .Q(out_slt_128), .SO(out_slt_128), .SE(scan_enable), .SI(out_slt_127));
SDFFNSRN u6_dout_reg_b8_b (.CK(clk_i), .D(n_11077), .Q(out_slt_129), .SO(out_slt_129), .SE(scan_enable), .SI(out_slt_128));
SDFFNSRN u6_dout_reg_b9_b (.CK(clk_i), .D(n_11076), .Q(out_slt_130), .SO(out_slt_130), .SE(scan_enable), .SI(out_slt_129));
SDFFNSRN u7_dout_reg_b10_b (.CK(clk_i), .D(n_11075), .Q(out_slt_150), .SO(out_slt_150), .SE(scan_enable), .SI(out_slt_130));
SDFFNSRN u7_dout_reg_b11_b (.CK(clk_i), .D(n_11074), .Q(out_slt_151), .SO(out_slt_151), .SE(scan_enable), .SI(out_slt_150));
SDFFNSRN u7_dout_reg_b12_b (.CK(clk_i), .D(n_11073), .Q(out_slt_152), .SO(out_slt_152), .SE(scan_enable), .SI(out_slt_151));
SDFFNSRN u7_dout_reg_b13_b (.CK(clk_i), .D(n_11072), .Q(out_slt_153), .SO(out_slt_153), .SE(scan_enable), .SI(out_slt_152));
SDFFNSRN u7_dout_reg_b14_b (.CK(clk_i), .D(n_11070), .Q(out_slt_154), .SO(out_slt_154), .SE(scan_enable), .SI(out_slt_153));
SDFFNSRN u7_dout_reg_b17_b (.CK(clk_i), .D(n_11065), .Q(out_slt_157), .SO(out_slt_157), .SE(scan_enable), .SI(out_slt_154));
SDFFNSRN u7_dout_reg_b15_b (.CK(clk_i), .D(n_11068), .Q(out_slt_155), .SO(out_slt_155), .SE(scan_enable), .SI(out_slt_157));
SDFFNSRN u7_dout_reg_b19_b (.CK(clk_i), .D(n_11063), .Q(out_slt_159), .SO(out_slt_159), .SE(scan_enable), .SI(out_slt_155));
SDFFNSRN u7_dout_reg_b16_b (.CK(clk_i), .D(n_11066), .Q(out_slt_156), .SO(out_slt_156), .SE(scan_enable), .SI(out_slt_159));
SDFFNSRN u7_dout_reg_b18_b (.CK(clk_i), .D(n_11064), .Q(out_slt_158), .SO(out_slt_158), .SE(scan_enable), .SI(out_slt_156));
SDFFNSRN u7_dout_reg_b4_b (.CK(clk_i), .D(n_11062), .Q(out_slt_144), .SO(out_slt_144), .SE(scan_enable), .SI(out_slt_158));
SDFFNSRN u7_dout_reg_b5_b (.CK(clk_i), .D(n_11061), .Q(out_slt_145), .SO(out_slt_145), .SE(scan_enable), .SI(out_slt_144));
SDFFNSRN u7_dout_reg_b6_b (.CK(clk_i), .D(n_11060), .Q(out_slt_146), .SO(out_slt_146), .SE(scan_enable), .SI(out_slt_145));
SDFFNSRN u7_dout_reg_b7_b (.CK(clk_i), .D(n_11058), .Q(out_slt_147), .SO(out_slt_147), .SE(scan_enable), .SI(out_slt_146));
SDFFNSRN u7_dout_reg_b8_b (.CK(clk_i), .D(n_11057), .Q(out_slt_148), .SO(out_slt_148), .SE(scan_enable), .SI(out_slt_147));
SDFFNSRN u7_dout_reg_b9_b (.CK(clk_i), .D(n_11056), .Q(out_slt_149), .SO(out_slt_149), .SE(scan_enable), .SI(out_slt_148));
SDFFNSRN u3_dout_reg_b10_b (.CK(clk_i), .D(n_11055), .Q(out_slt_74), .SO(out_slt_74), .SE(scan_enable), .SI(out_slt_149));
SDFFNSRN u3_dout_reg_b11_b (.CK(clk_i), .D(n_11054), .Q(out_slt_75), .SO(out_slt_75), .SE(scan_enable), .SI(out_slt_74));
SDFFNSRN u3_dout_reg_b13_b (.CK(clk_i), .D(n_11052), .Q(out_slt_77), .SO(out_slt_77), .SE(scan_enable), .SI(out_slt_75));
SDFFNSRN u3_dout_reg_b14_b (.CK(clk_i), .D(n_11051), .Q(out_slt_78), .SO(out_slt_78), .SE(scan_enable), .SI(out_slt_77));
SDFFNSRN u3_dout_reg_b15_b (.CK(clk_i), .D(n_11049), .Q(out_slt_79), .SO(out_slt_79), .SE(scan_enable), .SI(out_slt_78));
SDFFNSRN u3_dout_reg_b16_b (.CK(clk_i), .D(n_11047), .Q(out_slt_80), .SO(out_slt_80), .SE(scan_enable), .SI(out_slt_79));
SDFFNSRN u3_dout_reg_b17_b (.CK(clk_i), .D(n_11045), .Q(out_slt_81), .SO(out_slt_81), .SE(scan_enable), .SI(out_slt_80));
SDFFNSRN u3_dout_reg_b18_b (.CK(clk_i), .D(n_11044), .Q(out_slt_82), .SO(out_slt_82), .SE(scan_enable), .SI(out_slt_81));
SDFFNSRN u8_dout_reg_b10_b (.CK(clk_i), .D(n_11042), .Q(out_slt_169), .SO(out_slt_169), .SE(scan_enable), .SI(out_slt_82));
SDFFNSRN u3_dout_reg_b19_b (.CK(clk_i), .D(n_11041), .Q(out_slt_83), .SO(out_slt_83), .SE(scan_enable), .SI(out_slt_169));
SDFFNSRN u8_dout_reg_b11_b (.CK(clk_i), .D(n_11040), .Q(out_slt_170), .SO(out_slt_170), .SE(scan_enable), .SI(out_slt_83));
SDFFNSRN u8_dout_reg_b12_b (.CK(clk_i), .D(n_11039), .Q(out_slt_171), .SO(out_slt_171), .SE(scan_enable), .SI(out_slt_170));
SDFFNSRN u3_dout_reg_b12_b (.CK(clk_i), .D(n_11053), .Q(out_slt_76), .SO(out_slt_76), .SE(scan_enable), .SI(out_slt_171));
SDFFNSRN u8_dout_reg_b13_b (.CK(clk_i), .D(n_11038), .Q(out_slt_172), .SO(out_slt_172), .SE(scan_enable), .SI(out_slt_76));
SDFFNSRN u8_dout_reg_b14_b (.CK(clk_i), .D(n_11037), .Q(out_slt_173), .SO(out_slt_173), .SE(scan_enable), .SI(out_slt_172));
SDFFNSRN u3_dout_reg_b4_b (.CK(clk_i), .D(n_11035), .Q(out_slt_68), .SO(out_slt_68), .SE(scan_enable), .SI(out_slt_173));
SDFFNSRN u8_dout_reg_b16_b (.CK(clk_i), .D(n_11031), .Q(out_slt_175), .SO(out_slt_175), .SE(scan_enable), .SI(out_slt_68));
SDFFNSRN u3_dout_reg_b6_b (.CK(clk_i), .D(n_11028), .Q(out_slt_70), .SO(out_slt_70), .SE(scan_enable), .SI(out_slt_175));
SDFFNSRN u8_dout_reg_b17_b (.CK(clk_i), .D(n_11029), .Q(out_slt_176), .SO(out_slt_176), .SE(scan_enable), .SI(out_slt_70));
SDFFNSRN u3_dout_reg_b7_b (.CK(clk_i), .D(n_11027), .Q(out_slt_71), .SO(out_slt_71), .SE(scan_enable), .SI(out_slt_176));
SDFFNSRN u8_dout_reg_b18_b (.CK(clk_i), .D(n_11026), .Q(out_slt_177), .SO(out_slt_177), .SE(scan_enable), .SI(out_slt_71));
SDFFNSRN u3_dout_reg_b8_b (.CK(clk_i), .D(n_11024), .Q(out_slt_72), .SO(out_slt_72), .SE(scan_enable), .SI(out_slt_177));
SDFFNSRN u8_dout_reg_b15_b (.CK(clk_i), .D(n_11034), .Q(out_slt_174), .SO(out_slt_174), .SE(scan_enable), .SI(out_slt_72));
SDFFNSRN u3_dout_reg_b5_b (.CK(clk_i), .D(n_11032), .Q(out_slt_69), .SO(out_slt_69), .SE(scan_enable), .SI(out_slt_174));
SDFFNSRN u8_dout_reg_b19_b (.CK(clk_i), .D(n_11023), .Q(out_slt_178), .SO(out_slt_178), .SE(scan_enable), .SI(out_slt_69));
SDFFNSRN u3_dout_reg_b9_b (.CK(clk_i), .D(n_11022), .Q(out_slt_73), .SO(out_slt_73), .SE(scan_enable), .SI(out_slt_178));
SDFFNSRN u8_dout_reg_b4_b (.CK(clk_i), .D(n_11021), .Q(out_slt_163), .SO(out_slt_163), .SE(scan_enable), .SI(out_slt_73));
SDFFNSRN u8_dout_reg_b5_b (.CK(clk_i), .D(n_11020), .Q(out_slt_164), .SO(out_slt_164), .SE(scan_enable), .SI(out_slt_163));
SDFFNSRN u8_dout_reg_b6_b (.CK(clk_i), .D(n_11019), .Q(out_slt_165), .SO(out_slt_165), .SE(scan_enable), .SI(out_slt_164));
SDFFNSRN u8_dout_reg_b7_b (.CK(clk_i), .D(n_11018), .Q(out_slt_166), .SO(out_slt_166), .SE(scan_enable), .SI(out_slt_165));
SDFFNSRN u8_dout_reg_b8_b (.CK(clk_i), .D(n_11017), .Q(out_slt_167), .SO(out_slt_167), .SE(scan_enable), .SI(out_slt_166));
SDFFNSRN u8_dout_reg_b9_b (.CK(clk_i), .D(n_11016), .Q(out_slt_168), .SO(out_slt_168), .SE(scan_enable), .SI(out_slt_167));
SDFFNSRN u16_u1_dma_req_r1_reg (.CK(clk_i), .D(n_11159), .Q(u16_u1_dma_req_r1), .SO(u16_u1_dma_req_r1), .SE(scan_enable), .SI(out_slt_168));
SDFFNSRN u16_u3_dma_req_r1_reg (.CK(clk_i), .D(n_11158), .Q(u16_u3_dma_req_r1), .SO(u16_u3_dma_req_r1), .SE(scan_enable), .SI(u16_u1_dma_req_r1));
SDFFN u16_u8_dma_req_reg (.CK(clk_i), .D(n_11906), .Q(dma_req_o_b8_b), .SO(dma_req_o_b8_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u16_u3_dma_req_r1));
SDFFNSRN u4_dout_reg_b3_b (.CK(clk_i), .D(n_10998), .Q(out_slt_86), .SO(out_slt_86), .SE(scan_enable), .SI(dma_req_o_b8_b));
SDFFNSRN u5_dout_reg_b3_b (.CK(clk_i), .D(n_10995), .Q(out_slt_105), .SO(out_slt_105), .SE(scan_enable), .SI(out_slt_86));
SDFFNSRN u5_dout_reg_b2_b (.CK(clk_i), .D(n_10996), .Q(out_slt_104), .SO(out_slt_104), .SE(scan_enable), .SI(out_slt_105));
SDFFNSRN u4_dout_reg_b2_b (.CK(clk_i), .D(n_10999), .Q(out_slt_85), .SO(out_slt_85), .SE(scan_enable), .SI(out_slt_104));
SDFFNSRN u16_u0_dma_req_r1_reg (.CK(clk_i), .D(n_11125), .Q(u16_u0_dma_req_r1), .SO(u16_u0_dma_req_r1), .SE(scan_enable), .SI(out_slt_85));
SDFFNSRN u16_u2_dma_req_r1_reg (.CK(clk_i), .D(n_11124), .Q(u16_u2_dma_req_r1), .SO(u16_u2_dma_req_r1), .SE(scan_enable), .SI(u16_u0_dma_req_r1));
SDFFNSRN u16_u4_dma_req_r1_reg (.CK(clk_i), .D(n_11123), .Q(u16_u4_dma_req_r1), .SO(u16_u4_dma_req_r1), .SE(scan_enable), .SI(u16_u2_dma_req_r1));
SDFFNSRN u16_u5_dma_req_r1_reg (.CK(clk_i), .D(n_11122), .Q(u16_u5_dma_req_r1), .SO(u16_u5_dma_req_r1), .SE(scan_enable), .SI(u16_u4_dma_req_r1));
SDFFNSRN u4_dout_reg_b4_b (.CK(clk_i), .D(n_10933), .Q(out_slt_87), .SO(out_slt_87), .SE(scan_enable), .SI(u16_u5_dma_req_r1));
SDFFNSRN u11_wp_reg_b3_b (.CK(clk_i), .D(n_10900), .Q(u11_wp_b3_b), .SO(u11_wp_b3_b), .SE(scan_enable), .SI(out_slt_87));
SDFFN u16_u6_dma_req_reg (.CK(clk_i), .D(n_12373), .Q(dma_req_o_b6_b), .SO(dma_req_o_b6_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u11_wp_b3_b));
SDFFN u16_u7_dma_req_reg (.CK(clk_i), .D(n_12378), .Q(dma_req_o_b7_b), .SO(dma_req_o_b7_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(dma_req_o_b6_b));
SDFFNSRN u5_dout_reg_b0_b (.CK(clk_i), .D(n_10952), .Q(out_slt6), .SO(out_slt6), .SE(scan_enable), .SI(dma_req_o_b7_b));
SDFFNSRN u5_dout_reg_b1_b (.CK(clk_i), .D(n_10951), .Q(out_slt_103), .SO(out_slt_103), .SE(scan_enable), .SI(out_slt6));
SDFFNSRN u4_dout_reg_b1_b (.CK(clk_i), .D(n_10955), .Q(out_slt_84), .SO(out_slt_84), .SE(scan_enable), .SI(out_slt_103));
SDFFNSRN u4_dout_reg_b0_b (.CK(clk_i), .D(n_10956), .Q(out_slt4), .SO(out_slt4), .SE(scan_enable), .SI(out_slt_84));
SDFFNSRN u4_rp_reg_b0_b (.CK(clk_i), .D(n_10807), .Q(u4_rp_b0_b), .SO(u4_rp_b0_b), .SE(scan_enable), .SI(out_slt4));
SDFFNSRN u5_rp_reg_b0_b (.CK(clk_i), .D(n_10806), .Q(n_6091), .SO(n_6091), .SE(scan_enable), .SI(u4_rp_b0_b));
SDFFNSRN u11_mem_reg_b0_b_b18_b (.CK(clk_i), .D(n_10899), .Q(u11_mem_b0_b_167), .SO(u11_mem_b0_b_167), .SE(scan_enable), .SI(n_6091));
SDFFNSRN u11_mem_reg_b0_b_b19_b (.CK(clk_i), .D(n_10898), .Q(u11_mem_b0_b_168), .SO(u11_mem_b0_b_168), .SE(scan_enable), .SI(u11_mem_b0_b_167));
SDFFNSRN u11_mem_reg_b1_b_b18_b (.CK(clk_i), .D(n_10897), .Q(u11_mem_b1_b_136), .SO(u11_mem_b1_b_136), .SE(scan_enable), .SI(u11_mem_b0_b_168));
SDFFNSRN u11_mem_reg_b1_b_b19_b (.CK(clk_i), .D(n_10896), .Q(u11_mem_b1_b_137), .SO(u11_mem_b1_b_137), .SE(scan_enable), .SI(u11_mem_b1_b_136));
SDFFNSRN u11_mem_reg_b1_b_b20_b (.CK(clk_i), .D(n_10895), .Q(u11_mem_b1_b_138), .SO(u11_mem_b1_b_138), .SE(scan_enable), .SI(u11_mem_b1_b_137));
SDFFNSRN u11_mem_reg_b1_b_b21_b (.CK(clk_i), .D(n_10894), .Q(u11_mem_b1_b_139), .SO(u11_mem_b1_b_139), .SE(scan_enable), .SI(u11_mem_b1_b_138));
SDFFNSRN u11_mem_reg_b1_b_b22_b (.CK(clk_i), .D(n_10893), .Q(u11_mem_b1_b_140), .SO(u11_mem_b1_b_140), .SE(scan_enable), .SI(u11_mem_b1_b_139));
SDFFNSRN u11_mem_reg_b1_b_b23_b (.CK(clk_i), .D(n_10892), .Q(u11_mem_b1_b_141), .SO(u11_mem_b1_b_141), .SE(scan_enable), .SI(u11_mem_b1_b_140));
SDFFNSRN u11_mem_reg_b1_b_b24_b (.CK(clk_i), .D(n_10890), .Q(u11_mem_b1_b_142), .SO(u11_mem_b1_b_142), .SE(scan_enable), .SI(u11_mem_b1_b_141));
SDFFNSRN u11_mem_reg_b1_b_b25_b (.CK(clk_i), .D(n_10888), .Q(u11_mem_b1_b_143), .SO(u11_mem_b1_b_143), .SE(scan_enable), .SI(u11_mem_b1_b_142));
SDFFNSRN u11_mem_reg_b1_b_b26_b (.CK(clk_i), .D(n_10886), .Q(u11_mem_b1_b_144), .SO(u11_mem_b1_b_144), .SE(scan_enable), .SI(u11_mem_b1_b_143));
SDFFNSRN u11_mem_reg_b1_b_b27_b (.CK(clk_i), .D(n_10885), .Q(u11_mem_b1_b_145), .SO(u11_mem_b1_b_145), .SE(scan_enable), .SI(u11_mem_b1_b_144));
SDFFNSRN u11_mem_reg_b1_b_b28_b (.CK(clk_i), .D(n_10884), .Q(u11_mem_b1_b_146), .SO(u11_mem_b1_b_146), .SE(scan_enable), .SI(u11_mem_b1_b_145));
SDFFNSRN u11_mem_reg_b1_b_b29_b (.CK(clk_i), .D(n_10882), .Q(u11_mem_b1_b_147), .SO(u11_mem_b1_b_147), .SE(scan_enable), .SI(u11_mem_b1_b_146));
SDFFNSRN u11_mem_reg_b1_b_b30_b (.CK(clk_i), .D(n_10881), .Q(u11_mem_b1_b_148), .SO(u11_mem_b1_b_148), .SE(scan_enable), .SI(u11_mem_b1_b_147));
SDFFNSRN u11_mem_reg_b1_b_b31_b (.CK(clk_i), .D(n_10879), .Q(u11_mem_b1_b_149), .SO(u11_mem_b1_b_149), .SE(scan_enable), .SI(u11_mem_b1_b_148));
SDFFNSRN u11_mem_reg_b2_b_b18_b (.CK(clk_i), .D(n_10877), .Q(u11_mem_b2_b_105), .SO(u11_mem_b2_b_105), .SE(scan_enable), .SI(u11_mem_b1_b_149));
SDFFNSRN u11_mem_reg_b2_b_b19_b (.CK(clk_i), .D(n_10876), .Q(u11_mem_b2_b_106), .SO(u11_mem_b2_b_106), .SE(scan_enable), .SI(u11_mem_b2_b_105));
SDFFNSRN u11_mem_reg_b2_b_b20_b (.CK(clk_i), .D(n_10875), .Q(u11_mem_b2_b_107), .SO(u11_mem_b2_b_107), .SE(scan_enable), .SI(u11_mem_b2_b_106));
SDFFNSRN u11_mem_reg_b2_b_b21_b (.CK(clk_i), .D(n_10873), .Q(u11_mem_b2_b_108), .SO(u11_mem_b2_b_108), .SE(scan_enable), .SI(u11_mem_b2_b_107));
SDFFNSRN u11_mem_reg_b2_b_b22_b (.CK(clk_i), .D(n_10872), .Q(u11_mem_b2_b_109), .SO(u11_mem_b2_b_109), .SE(scan_enable), .SI(u11_mem_b2_b_108));
SDFFNSRN u11_mem_reg_b2_b_b23_b (.CK(clk_i), .D(n_10870), .Q(u11_mem_b2_b_110), .SO(u11_mem_b2_b_110), .SE(scan_enable), .SI(u11_mem_b2_b_109));
SDFFNSRN u11_mem_reg_b2_b_b24_b (.CK(clk_i), .D(n_10868), .Q(u11_mem_b2_b_111), .SO(u11_mem_b2_b_111), .SE(scan_enable), .SI(u11_mem_b2_b_110));
SDFFNSRN u11_mem_reg_b2_b_b25_b (.CK(clk_i), .D(n_10867), .Q(u11_mem_b2_b_112), .SO(u11_mem_b2_b_112), .SE(scan_enable), .SI(u11_mem_b2_b_111));
SDFFNSRN u11_mem_reg_b2_b_b26_b (.CK(clk_i), .D(n_10866), .Q(u11_mem_b2_b_113), .SO(u11_mem_b2_b_113), .SE(scan_enable), .SI(u11_mem_b2_b_112));
SDFFNSRN u11_mem_reg_b2_b_b27_b (.CK(clk_i), .D(n_10864), .Q(u11_mem_b2_b_114), .SO(u11_mem_b2_b_114), .SE(scan_enable), .SI(u11_mem_b2_b_113));
SDFFNSRN u11_mem_reg_b2_b_b28_b (.CK(clk_i), .D(n_10863), .Q(u11_mem_b2_b_115), .SO(u11_mem_b2_b_115), .SE(scan_enable), .SI(u11_mem_b2_b_114));
SDFFNSRN u11_mem_reg_b2_b_b29_b (.CK(clk_i), .D(n_10862), .Q(u11_mem_b2_b_116), .SO(u11_mem_b2_b_116), .SE(scan_enable), .SI(u11_mem_b2_b_115));
SDFFNSRN u11_mem_reg_b2_b_b30_b (.CK(clk_i), .D(n_10860), .Q(u11_mem_b2_b_117), .SO(u11_mem_b2_b_117), .SE(scan_enable), .SI(u11_mem_b2_b_116));
SDFFNSRN u11_mem_reg_b2_b_b31_b (.CK(clk_i), .D(n_10859), .Q(u11_mem_b2_b_118), .SO(u11_mem_b2_b_118), .SE(scan_enable), .SI(u11_mem_b2_b_117));
SDFFNSRN u11_mem_reg_b3_b_b18_b (.CK(clk_i), .D(n_10858), .Q(u11_mem_b3_b_74), .SO(u11_mem_b3_b_74), .SE(scan_enable), .SI(u11_mem_b2_b_118));
SDFFNSRN u11_mem_reg_b3_b_b19_b (.CK(clk_i), .D(n_10857), .Q(u11_mem_b3_b_75), .SO(u11_mem_b3_b_75), .SE(scan_enable), .SI(u11_mem_b3_b_74));
SDFFNSRN u11_mem_reg_b3_b_b20_b (.CK(clk_i), .D(n_10856), .Q(u11_mem_b3_b_76), .SO(u11_mem_b3_b_76), .SE(scan_enable), .SI(u11_mem_b3_b_75));
SDFFNSRN u11_mem_reg_b3_b_b21_b (.CK(clk_i), .D(n_10855), .Q(u11_mem_b3_b_77), .SO(u11_mem_b3_b_77), .SE(scan_enable), .SI(u11_mem_b3_b_76));
SDFFNSRN u11_mem_reg_b3_b_b22_b (.CK(clk_i), .D(n_10854), .Q(u11_mem_b3_b_78), .SO(u11_mem_b3_b_78), .SE(scan_enable), .SI(u11_mem_b3_b_77));
SDFFNSRN u11_mem_reg_b3_b_b23_b (.CK(clk_i), .D(n_10853), .Q(u11_mem_b3_b_79), .SO(u11_mem_b3_b_79), .SE(scan_enable), .SI(u11_mem_b3_b_78));
SDFFNSRN u11_mem_reg_b3_b_b24_b (.CK(clk_i), .D(n_10852), .Q(u11_mem_b3_b_80), .SO(u11_mem_b3_b_80), .SE(scan_enable), .SI(u11_mem_b3_b_79));
SDFFNSRN u11_mem_reg_b3_b_b25_b (.CK(clk_i), .D(n_10851), .Q(u11_mem_b3_b_81), .SO(u11_mem_b3_b_81), .SE(scan_enable), .SI(u11_mem_b3_b_80));
SDFFNSRN u11_mem_reg_b3_b_b26_b (.CK(clk_i), .D(n_10850), .Q(u11_mem_b3_b_82), .SO(u11_mem_b3_b_82), .SE(scan_enable), .SI(u11_mem_b3_b_81));
SDFFNSRN u11_mem_reg_b3_b_b27_b (.CK(clk_i), .D(n_10849), .Q(u11_mem_b3_b_83), .SO(u11_mem_b3_b_83), .SE(scan_enable), .SI(u11_mem_b3_b_82));
SDFFNSRN u11_mem_reg_b3_b_b28_b (.CK(clk_i), .D(n_10848), .Q(u11_mem_b3_b_84), .SO(u11_mem_b3_b_84), .SE(scan_enable), .SI(u11_mem_b3_b_83));
SDFFNSRN u11_mem_reg_b3_b_b29_b (.CK(clk_i), .D(n_10847), .Q(u11_mem_b3_b_85), .SO(u11_mem_b3_b_85), .SE(scan_enable), .SI(u11_mem_b3_b_84));
SDFFNSRN u11_mem_reg_b3_b_b30_b (.CK(clk_i), .D(n_10846), .Q(u11_mem_b3_b_86), .SO(u11_mem_b3_b_86), .SE(scan_enable), .SI(u11_mem_b3_b_85));
SDFFNSRN u11_mem_reg_b3_b_b31_b (.CK(clk_i), .D(n_10845), .Q(u11_mem_b3_b_87), .SO(u11_mem_b3_b_87), .SE(scan_enable), .SI(u11_mem_b3_b_86));
SDFFNSRN u11_mem_reg_b3_b_b7_b (.CK(clk_i), .D(n_10827), .Q(u11_mem_b3_b_63), .SO(u11_mem_b3_b_63), .SE(scan_enable), .SI(u11_mem_b3_b_87));
SDFFNSRN u11_mem_reg_b1_b_b12_b (.CK(clk_i), .D(n_10844), .Q(u11_mem_b1_b_130), .SO(u11_mem_b1_b_130), .SE(scan_enable), .SI(u11_mem_b3_b_63));
SDFFNSRN u11_mem_reg_b1_b_b13_b (.CK(clk_i), .D(n_10843), .Q(u11_mem_b1_b_131), .SO(u11_mem_b1_b_131), .SE(scan_enable), .SI(u11_mem_b1_b_130));
SDFFNSRN u11_mem_reg_b1_b_b16_b (.CK(clk_i), .D(n_10842), .Q(u11_mem_b1_b_134), .SO(u11_mem_b1_b_134), .SE(scan_enable), .SI(u11_mem_b1_b_131));
SDFFNSRN u11_mem_reg_b2_b_b17_b (.CK(clk_i), .D(n_10841), .Q(u11_mem_b2_b_104), .SO(u11_mem_b2_b_104), .SE(scan_enable), .SI(u11_mem_b1_b_134));
SDFFNSRN u11_mem_reg_b2_b_b1_b (.CK(clk_i), .D(n_10840), .Q(u11_mem_b2_b_88), .SO(u11_mem_b2_b_88), .SE(scan_enable), .SI(u11_mem_b2_b_104));
SDFFNSRN u11_mem_reg_b2_b_b7_b (.CK(clk_i), .D(n_10838), .Q(u11_mem_b2_b_94), .SO(u11_mem_b2_b_94), .SE(scan_enable), .SI(u11_mem_b2_b_88));
SDFFNSRN u11_mem_reg_b2_b_b8_b (.CK(clk_i), .D(n_10837), .Q(u11_mem_b2_b_95), .SO(u11_mem_b2_b_95), .SE(scan_enable), .SI(u11_mem_b2_b_94));
SDFFNSRN u11_mem_reg_b3_b_b16_b (.CK(clk_i), .D(n_10836), .Q(u11_mem_b3_b_72), .SO(u11_mem_b3_b_72), .SE(scan_enable), .SI(u11_mem_b2_b_95));
SDFFNSRN u11_mem_reg_b3_b_b17_b (.CK(clk_i), .D(n_10834), .Q(u11_mem_b3_b_73), .SO(u11_mem_b3_b_73), .SE(scan_enable), .SI(u11_mem_b3_b_72));
SDFFNSRN u11_mem_reg_b3_b_b5_b (.CK(clk_i), .D(n_10829), .Q(u11_mem_b3_b_61), .SO(u11_mem_b3_b_61), .SE(scan_enable), .SI(u11_mem_b3_b_73));
SDFFNSRN u11_mem_reg_b3_b_b6_b (.CK(clk_i), .D(n_10828), .Q(u11_mem_b3_b_62), .SO(u11_mem_b3_b_62), .SE(scan_enable), .SI(u11_mem_b3_b_61));
SDFFNSRN u11_wp_reg_b1_b (.CK(clk_i), .D(n_10902), .Q(u11_wp_b1_b), .SO(u11_wp_b1_b), .SE(scan_enable), .SI(u11_mem_b3_b_62));
SDFFNSRN u11_wp_reg_b2_b (.CK(clk_i), .D(n_10948), .Q(u11_wp_b2_b), .SO(u11_wp_b2_b), .SE(scan_enable), .SI(u11_wp_b1_b));
SDFFNSRN u4_dout_reg_b10_b (.CK(clk_i), .D(n_10947), .Q(out_slt_93), .SO(out_slt_93), .SE(scan_enable), .SI(u11_wp_b2_b));
SDFFNSRN u4_dout_reg_b13_b (.CK(clk_i), .D(n_10943), .Q(out_slt_96), .SO(out_slt_96), .SE(scan_enable), .SI(out_slt_93));
SDFFNSRN u4_dout_reg_b14_b (.CK(clk_i), .D(n_10942), .Q(out_slt_97), .SO(out_slt_97), .SE(scan_enable), .SI(out_slt_96));
SDFFNSRN u4_dout_reg_b15_b (.CK(clk_i), .D(n_10941), .Q(out_slt_98), .SO(out_slt_98), .SE(scan_enable), .SI(out_slt_97));
SDFFNSRN u4_dout_reg_b16_b (.CK(clk_i), .D(n_10939), .Q(out_slt_99), .SO(out_slt_99), .SE(scan_enable), .SI(out_slt_98));
SDFFNSRN u4_dout_reg_b11_b (.CK(clk_i), .D(n_10946), .Q(out_slt_94), .SO(out_slt_94), .SE(scan_enable), .SI(out_slt_99));
SDFFNSRN u4_dout_reg_b18_b (.CK(clk_i), .D(n_10935), .Q(out_slt_101), .SO(out_slt_101), .SE(scan_enable), .SI(out_slt_94));
SDFFNSRN u4_dout_reg_b12_b (.CK(clk_i), .D(n_10944), .Q(out_slt_95), .SO(out_slt_95), .SE(scan_enable), .SI(out_slt_101));
SDFFNSRN u4_dout_reg_b19_b (.CK(clk_i), .D(n_10934), .Q(out_slt_102), .SO(out_slt_102), .SE(scan_enable), .SI(out_slt_95));
SDFFNSRN u4_dout_reg_b17_b (.CK(clk_i), .D(n_10937), .Q(out_slt_100), .SO(out_slt_100), .SE(scan_enable), .SI(out_slt_102));
SDFFNSRN u4_dout_reg_b5_b (.CK(clk_i), .D(n_10932), .Q(out_slt_88), .SO(out_slt_88), .SE(scan_enable), .SI(out_slt_100));
SDFFNSRN u4_dout_reg_b6_b (.CK(clk_i), .D(n_10931), .Q(out_slt_89), .SO(out_slt_89), .SE(scan_enable), .SI(out_slt_88));
SDFFNSRN u4_dout_reg_b7_b (.CK(clk_i), .D(n_10930), .Q(out_slt_90), .SO(out_slt_90), .SE(scan_enable), .SI(out_slt_89));
SDFFNSRN u4_dout_reg_b8_b (.CK(clk_i), .D(n_10929), .Q(out_slt_91), .SO(out_slt_91), .SE(scan_enable), .SI(out_slt_90));
SDFFNSRN u4_dout_reg_b9_b (.CK(clk_i), .D(n_10928), .Q(out_slt_92), .SO(out_slt_92), .SE(scan_enable), .SI(out_slt_91));
SDFFNSRN u5_dout_reg_b10_b (.CK(clk_i), .D(n_10927), .Q(out_slt_112), .SO(out_slt_112), .SE(scan_enable), .SI(out_slt_92));
SDFFNSRN u5_dout_reg_b11_b (.CK(clk_i), .D(n_10926), .Q(out_slt_113), .SO(out_slt_113), .SE(scan_enable), .SI(out_slt_112));
SDFFNSRN u5_dout_reg_b12_b (.CK(clk_i), .D(n_10924), .Q(out_slt_114), .SO(out_slt_114), .SE(scan_enable), .SI(out_slt_113));
SDFFNSRN u5_dout_reg_b14_b (.CK(clk_i), .D(n_10922), .Q(out_slt_116), .SO(out_slt_116), .SE(scan_enable), .SI(out_slt_114));
SDFFNSRN u5_dout_reg_b15_b (.CK(clk_i), .D(n_10920), .Q(out_slt_117), .SO(out_slt_117), .SE(scan_enable), .SI(out_slt_116));
SDFFNSRN u5_dout_reg_b16_b (.CK(clk_i), .D(n_10919), .Q(out_slt_118), .SO(out_slt_118), .SE(scan_enable), .SI(out_slt_117));
SDFFNSRN u5_dout_reg_b18_b (.CK(clk_i), .D(n_10915), .Q(out_slt_120), .SO(out_slt_120), .SE(scan_enable), .SI(out_slt_118));
SDFFNSRN u5_dout_reg_b19_b (.CK(clk_i), .D(n_10914), .Q(out_slt_121), .SO(out_slt_121), .SE(scan_enable), .SI(out_slt_120));
SDFFNSRN u5_dout_reg_b4_b (.CK(clk_i), .D(n_10913), .Q(out_slt_106), .SO(out_slt_106), .SE(scan_enable), .SI(out_slt_121));
SDFFNSRN u5_dout_reg_b5_b (.CK(clk_i), .D(n_10912), .Q(out_slt_107), .SO(out_slt_107), .SE(scan_enable), .SI(out_slt_106));
SDFFNSRN u5_dout_reg_b6_b (.CK(clk_i), .D(n_10911), .Q(out_slt_108), .SO(out_slt_108), .SE(scan_enable), .SI(out_slt_107));
SDFFNSRN u5_dout_reg_b8_b (.CK(clk_i), .D(n_10909), .Q(out_slt_110), .SO(out_slt_110), .SE(scan_enable), .SI(out_slt_108));
SDFFNSRN u5_dout_reg_b9_b (.CK(clk_i), .D(n_10908), .Q(out_slt_111), .SO(out_slt_111), .SE(scan_enable), .SI(out_slt_110));
SDFFNSRN u11_mem_reg_b0_b_b0_b (.CK(clk_i), .D(n_10821), .Q(u11_mem_b0_b), .SO(u11_mem_b0_b), .SE(scan_enable), .SI(out_slt_111));
SDFFNSRN u11_mem_reg_b0_b_b10_b (.CK(clk_i), .D(n_10819), .Q(u11_mem_b0_b_159), .SO(u11_mem_b0_b_159), .SE(scan_enable), .SI(u11_mem_b0_b));
SDFFNSRN u11_mem_reg_b0_b_b11_b (.CK(clk_i), .D(n_10818), .Q(u11_mem_b0_b_160), .SO(u11_mem_b0_b_160), .SE(scan_enable), .SI(u11_mem_b0_b_159));
SDFFNSRN u11_mem_reg_b0_b_b12_b (.CK(clk_i), .D(n_10815), .Q(u11_mem_b0_b_161), .SO(u11_mem_b0_b_161), .SE(scan_enable), .SI(u11_mem_b0_b_160));
SDFFNSRN u11_mem_reg_b0_b_b13_b (.CK(clk_i), .D(n_10817), .Q(u11_mem_b0_b_162), .SO(u11_mem_b0_b_162), .SE(scan_enable), .SI(u11_mem_b0_b_161));
SDFFNSRN u11_mem_reg_b0_b_b14_b (.CK(clk_i), .D(n_10814), .Q(u11_mem_b0_b_163), .SO(u11_mem_b0_b_163), .SE(scan_enable), .SI(u11_mem_b0_b_162));
SDFFNSRN u11_mem_reg_b0_b_b15_b (.CK(clk_i), .D(n_10813), .Q(u11_mem_b0_b_164), .SO(u11_mem_b0_b_164), .SE(scan_enable), .SI(u11_mem_b0_b_163));
SDFFNSRN u11_mem_reg_b0_b_b1_b (.CK(clk_i), .D(n_10812), .Q(u11_mem_b0_b_150), .SO(u11_mem_b0_b_150), .SE(scan_enable), .SI(u11_mem_b0_b_164));
SDFFN u15_crac_rd_reg (.CK(clk_i), .D(n_10903), .Q(u15_crac_rd), .SO(u15_crac_rd), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u11_mem_b0_b_150));
SDFFN u17_int_set_reg_b1_b (.CK(clk_i), .D(n_10907), .Q(oc0_int_set_707), .SO(oc0_int_set_707), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u15_crac_rd));
SDFFN u20_int_set_reg_b1_b (.CK(clk_i), .D(n_10906), .Q(oc3_int_set_713), .SO(oc3_int_set_713), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc0_int_set_707));
SDFFN u21_int_set_reg_b1_b (.CK(clk_i), .D(n_10905), .Q(oc4_int_set_715), .SO(oc4_int_set_715), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc3_int_set_713));
SDFFN u22_int_set_reg_b1_b (.CK(clk_i), .D(n_10904), .Q(oc5_int_set_717), .SO(oc5_int_set_717), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc4_int_set_715));
SDFFNSRN u5_dout_reg_b7_b (.CK(clk_i), .D(n_10910), .Q(out_slt_109), .SO(out_slt_109), .SE(scan_enable), .SI(oc5_int_set_717));
SDFFNSRN u5_dout_reg_b17_b (.CK(clk_i), .D(n_10917), .Q(out_slt_119), .SO(out_slt_119), .SE(scan_enable), .SI(out_slt_109));
SDFFNSRN u5_dout_reg_b13_b (.CK(clk_i), .D(n_10923), .Q(out_slt_115), .SO(out_slt_115), .SE(scan_enable), .SI(out_slt_119));
SDFFNSRN u10_mem_reg_b0_b_b18_b (.CK(clk_i), .D(n_10678), .Q(u10_mem_b0_b_167), .SO(u10_mem_b0_b_167), .SE(scan_enable), .SI(out_slt_115));
SDFFNSRN u10_mem_reg_b3_b_b28_b (.CK(clk_i), .D(n_10684), .Q(u10_mem_b3_b_84), .SO(u10_mem_b3_b_84), .SE(scan_enable), .SI(u10_mem_b0_b_167));
SDFFNSRN u10_mem_reg_b3_b_b24_b (.CK(clk_i), .D(n_10690), .Q(u10_mem_b3_b_80), .SO(u10_mem_b3_b_80), .SE(scan_enable), .SI(u10_mem_b3_b_84));
SDFFNSRN u9_mem_reg_b3_b_b30_b (.CK(clk_i), .D(n_10701), .Q(u9_mem_b3_b_86), .SO(u9_mem_b3_b_86), .SE(scan_enable), .SI(u10_mem_b3_b_80));
SDFFNSRN u9_mem_reg_b3_b_b26_b (.CK(clk_i), .D(n_10705), .Q(u9_mem_b3_b_82), .SO(u9_mem_b3_b_82), .SE(scan_enable), .SI(u9_mem_b3_b_86));
SDFFNSRN u10_wp_reg_b3_b (.CK(clk_i), .D(n_10778), .Q(u10_wp_b3_b), .SO(u10_wp_b3_b), .SE(scan_enable), .SI(u9_mem_b3_b_82));
SDFFNSRN u9_mem_reg_b3_b_b22_b (.CK(clk_i), .D(n_10709), .Q(u9_mem_b3_b_78), .SO(u9_mem_b3_b_78), .SE(scan_enable), .SI(u10_wp_b3_b));
SDFFNSRN u9_mem_reg_b2_b_b28_b (.CK(clk_i), .D(n_10718), .Q(u9_mem_b2_b_115), .SO(u9_mem_b2_b_115), .SE(scan_enable), .SI(u9_mem_b3_b_78));
SDFFNSRN u9_mem_reg_b2_b_b24_b (.CK(clk_i), .D(n_10723), .Q(u9_mem_b2_b_111), .SO(u9_mem_b2_b_111), .SE(scan_enable), .SI(u9_mem_b2_b_115));
SDFFNSRN u9_mem_reg_b2_b_b20_b (.CK(clk_i), .D(n_10730), .Q(u9_mem_b2_b_107), .SO(u9_mem_b2_b_107), .SE(scan_enable), .SI(u9_mem_b2_b_111));
SDFFNSRN u9_mem_reg_b1_b_b28_b (.CK(clk_i), .D(n_10742), .Q(u9_mem_b1_b_146), .SO(u9_mem_b1_b_146), .SE(scan_enable), .SI(u9_mem_b2_b_107));
SDFFNSRN u9_mem_reg_b1_b_b25_b (.CK(clk_i), .D(n_10746), .Q(u9_mem_b1_b_143), .SO(u9_mem_b1_b_143), .SE(scan_enable), .SI(u9_mem_b1_b_146));
SDFFNSRN u9_mem_reg_b1_b_b22_b (.CK(clk_i), .D(n_10751), .Q(u9_mem_b1_b_140), .SO(u9_mem_b1_b_140), .SE(scan_enable), .SI(u9_mem_b1_b_143));
SDFFNSRN u10_mem_reg_b2_b_b24_b (.CK(clk_i), .D(n_10763), .Q(u10_mem_b2_b_111), .SO(u10_mem_b2_b_111), .SE(scan_enable), .SI(u9_mem_b1_b_140));
SDFFNSRN u11_mem_reg_b3_b_b14_b (.CK(clk_i), .D(n_10457), .Q(u11_mem_b3_b_70), .SO(u11_mem_b3_b_70), .SE(scan_enable), .SI(u10_mem_b2_b_111));
SDFFNSRN u11_mem_reg_b3_b_b0_b (.CK(clk_i), .D(n_10472), .Q(u11_mem_b3_b), .SO(u11_mem_b3_b), .SE(scan_enable), .SI(u11_mem_b3_b_70));
SDFFNSRN u11_mem_reg_b3_b_b13_b (.CK(clk_i), .D(n_10458), .Q(u11_mem_b3_b_69), .SO(u11_mem_b3_b_69), .SE(scan_enable), .SI(u11_mem_b3_b));
SDFFNSRN u10_mem_reg_b1_b_b0_b (.CK(clk_i), .D(n_10544), .Q(u10_mem_b1_b), .SO(u10_mem_b1_b), .SE(scan_enable), .SI(u11_mem_b3_b_69));
SDFFNSRN u11_mem_reg_b1_b_b15_b (.CK(clk_i), .D(n_10558), .Q(u11_mem_b1_b_133), .SO(u11_mem_b1_b_133), .SE(scan_enable), .SI(u10_mem_b1_b));
SDFFNSRN u11_mem_reg_b1_b_b6_b (.CK(clk_i), .D(n_10547), .Q(u11_mem_b1_b_124), .SO(u11_mem_b1_b_124), .SE(scan_enable), .SI(u11_mem_b1_b_133));
SDFFNSRN u10_mem_reg_b2_b_b18_b (.CK(clk_i), .D(n_10772), .Q(u10_mem_b2_b_105), .SO(u10_mem_b2_b_105), .SE(scan_enable), .SI(u11_mem_b1_b_124));
SDFFNSRN u10_mem_reg_b2_b_b19_b (.CK(clk_i), .D(n_10771), .Q(u10_mem_b2_b_106), .SO(u10_mem_b2_b_106), .SE(scan_enable), .SI(u10_mem_b2_b_105));
SDFFNSRN u10_mem_reg_b2_b_b20_b (.CK(clk_i), .D(n_10770), .Q(u10_mem_b2_b_107), .SO(u10_mem_b2_b_107), .SE(scan_enable), .SI(u10_mem_b2_b_106));
SDFFNSRN u10_mem_reg_b2_b_b21_b (.CK(clk_i), .D(n_10769), .Q(u10_mem_b2_b_108), .SO(u10_mem_b2_b_108), .SE(scan_enable), .SI(u10_mem_b2_b_107));
SDFFNSRN u10_mem_reg_b2_b_b22_b (.CK(clk_i), .D(n_10768), .Q(u10_mem_b2_b_109), .SO(u10_mem_b2_b_109), .SE(scan_enable), .SI(u10_mem_b2_b_108));
SDFFNSRN u9_mem_reg_b0_b_b18_b (.CK(clk_i), .D(n_10765), .Q(u9_mem_b0_b_167), .SO(u9_mem_b0_b_167), .SE(scan_enable), .SI(u10_mem_b2_b_109));
SDFFNSRN u9_mem_reg_b0_b_b19_b (.CK(clk_i), .D(n_10764), .Q(u9_mem_b0_b_168), .SO(u9_mem_b0_b_168), .SE(scan_enable), .SI(u9_mem_b0_b_167));
SDFFNSRN u10_mem_reg_b2_b_b23_b (.CK(clk_i), .D(n_10766), .Q(u10_mem_b2_b_110), .SO(u10_mem_b2_b_110), .SE(scan_enable), .SI(u9_mem_b0_b_168));
SDFFNSRN u10_mem_reg_b2_b_b25_b (.CK(clk_i), .D(n_10762), .Q(u10_mem_b2_b_112), .SO(u10_mem_b2_b_112), .SE(scan_enable), .SI(u10_mem_b2_b_110));
SDFFNSRN u10_mem_reg_b2_b_b26_b (.CK(clk_i), .D(n_10760), .Q(u10_mem_b2_b_113), .SO(u10_mem_b2_b_113), .SE(scan_enable), .SI(u10_mem_b2_b_112));
SDFFNSRN u10_mem_reg_b2_b_b27_b (.CK(clk_i), .D(n_10758), .Q(u10_mem_b2_b_114), .SO(u10_mem_b2_b_114), .SE(scan_enable), .SI(u10_mem_b2_b_113));
SDFFNSRN u9_mem_reg_b1_b_b18_b (.CK(clk_i), .D(n_10756), .Q(u9_mem_b1_b_136), .SO(u9_mem_b1_b_136), .SE(scan_enable), .SI(u10_mem_b2_b_114));
SDFFNSRN u9_mem_reg_b1_b_b19_b (.CK(clk_i), .D(n_10755), .Q(u9_mem_b1_b_137), .SO(u9_mem_b1_b_137), .SE(scan_enable), .SI(u9_mem_b1_b_136));
SDFFNSRN u9_mem_reg_b1_b_b20_b (.CK(clk_i), .D(n_10754), .Q(u9_mem_b1_b_138), .SO(u9_mem_b1_b_138), .SE(scan_enable), .SI(u9_mem_b1_b_137));
SDFFNSRN u9_mem_reg_b1_b_b21_b (.CK(clk_i), .D(n_10753), .Q(u9_mem_b1_b_139), .SO(u9_mem_b1_b_139), .SE(scan_enable), .SI(u9_mem_b1_b_138));
SDFFNSRN u10_mem_reg_b2_b_b28_b (.CK(clk_i), .D(n_10757), .Q(u10_mem_b2_b_115), .SO(u10_mem_b2_b_115), .SE(scan_enable), .SI(u9_mem_b1_b_139));
SDFFNSRN u9_mem_reg_b1_b_b23_b (.CK(clk_i), .D(n_10750), .Q(u9_mem_b1_b_141), .SO(u9_mem_b1_b_141), .SE(scan_enable), .SI(u10_mem_b2_b_115));
SDFFNSRN u9_mem_reg_b1_b_b24_b (.CK(clk_i), .D(n_10748), .Q(u9_mem_b1_b_142), .SO(u9_mem_b1_b_142), .SE(scan_enable), .SI(u9_mem_b1_b_141));
SDFFNSRN u9_mem_reg_b1_b_b26_b (.CK(clk_i), .D(n_10744), .Q(u9_mem_b1_b_144), .SO(u9_mem_b1_b_144), .SE(scan_enable), .SI(u9_mem_b1_b_142));
SDFFNSRN u10_mem_reg_b2_b_b29_b (.CK(clk_i), .D(n_10752), .Q(u10_mem_b2_b_116), .SO(u10_mem_b2_b_116), .SE(scan_enable), .SI(u9_mem_b1_b_144));
SDFFNSRN u9_mem_reg_b1_b_b27_b (.CK(clk_i), .D(n_10743), .Q(u9_mem_b1_b_145), .SO(u9_mem_b1_b_145), .SE(scan_enable), .SI(u10_mem_b2_b_116));
SDFFNSRN u9_mem_reg_b1_b_b29_b (.CK(clk_i), .D(n_10740), .Q(u9_mem_b1_b_147), .SO(u9_mem_b1_b_147), .SE(scan_enable), .SI(u9_mem_b1_b_145));
SDFFNSRN u9_mem_reg_b1_b_b30_b (.CK(clk_i), .D(n_10739), .Q(u9_mem_b1_b_148), .SO(u9_mem_b1_b_148), .SE(scan_enable), .SI(u9_mem_b1_b_147));
SDFFNSRN u9_mem_reg_b1_b_b31_b (.CK(clk_i), .D(n_10737), .Q(u9_mem_b1_b_149), .SO(u9_mem_b1_b_149), .SE(scan_enable), .SI(u9_mem_b1_b_148));
SDFFNSRN u10_mem_reg_b2_b_b30_b (.CK(clk_i), .D(n_10735), .Q(u10_mem_b2_b_117), .SO(u10_mem_b2_b_117), .SE(scan_enable), .SI(u9_mem_b1_b_149));
SDFFNSRN u9_mem_reg_b2_b_b18_b (.CK(clk_i), .D(n_10732), .Q(u9_mem_b2_b_105), .SO(u9_mem_b2_b_105), .SE(scan_enable), .SI(u10_mem_b2_b_117));
SDFFNSRN u9_mem_reg_b2_b_b19_b (.CK(clk_i), .D(n_10731), .Q(u9_mem_b2_b_106), .SO(u9_mem_b2_b_106), .SE(scan_enable), .SI(u9_mem_b2_b_105));
SDFFNSRN u10_mem_reg_b2_b_b31_b (.CK(clk_i), .D(n_10733), .Q(u10_mem_b2_b_118), .SO(u10_mem_b2_b_118), .SE(scan_enable), .SI(u9_mem_b2_b_106));
SDFFNSRN u9_mem_reg_b2_b_b21_b (.CK(clk_i), .D(n_10728), .Q(u9_mem_b2_b_108), .SO(u9_mem_b2_b_108), .SE(scan_enable), .SI(u10_mem_b2_b_118));
SDFFNSRN u9_mem_reg_b2_b_b22_b (.CK(clk_i), .D(n_10727), .Q(u9_mem_b2_b_109), .SO(u9_mem_b2_b_109), .SE(scan_enable), .SI(u9_mem_b2_b_108));
SDFFNSRN u9_mem_reg_b2_b_b23_b (.CK(clk_i), .D(n_10725), .Q(u9_mem_b2_b_110), .SO(u9_mem_b2_b_110), .SE(scan_enable), .SI(u9_mem_b2_b_109));
SDFFNSRN u9_mem_reg_b2_b_b25_b (.CK(clk_i), .D(n_10722), .Q(u9_mem_b2_b_112), .SO(u9_mem_b2_b_112), .SE(scan_enable), .SI(u9_mem_b2_b_110));
SDFFNSRN u9_mem_reg_b2_b_b26_b (.CK(clk_i), .D(n_10721), .Q(u9_mem_b2_b_113), .SO(u9_mem_b2_b_113), .SE(scan_enable), .SI(u9_mem_b2_b_112));
SDFFNSRN u9_mem_reg_b2_b_b27_b (.CK(clk_i), .D(n_10719), .Q(u9_mem_b2_b_114), .SO(u9_mem_b2_b_114), .SE(scan_enable), .SI(u9_mem_b2_b_113));
SDFFNSRN u9_mem_reg_b2_b_b29_b (.CK(clk_i), .D(n_10717), .Q(u9_mem_b2_b_116), .SO(u9_mem_b2_b_116), .SE(scan_enable), .SI(u9_mem_b2_b_114));
SDFFNSRN u9_mem_reg_b2_b_b30_b (.CK(clk_i), .D(n_10715), .Q(u9_mem_b2_b_117), .SO(u9_mem_b2_b_117), .SE(scan_enable), .SI(u9_mem_b2_b_116));
SDFFNSRN u9_mem_reg_b2_b_b31_b (.CK(clk_i), .D(n_10714), .Q(u9_mem_b2_b_118), .SO(u9_mem_b2_b_118), .SE(scan_enable), .SI(u9_mem_b2_b_117));
SDFFNSRN u9_mem_reg_b3_b_b18_b (.CK(clk_i), .D(n_10713), .Q(u9_mem_b3_b_74), .SO(u9_mem_b3_b_74), .SE(scan_enable), .SI(u9_mem_b2_b_118));
SDFFNSRN u9_mem_reg_b3_b_b19_b (.CK(clk_i), .D(n_10712), .Q(u9_mem_b3_b_75), .SO(u9_mem_b3_b_75), .SE(scan_enable), .SI(u9_mem_b3_b_74));
SDFFNSRN u9_mem_reg_b3_b_b20_b (.CK(clk_i), .D(n_10711), .Q(u9_mem_b3_b_76), .SO(u9_mem_b3_b_76), .SE(scan_enable), .SI(u9_mem_b3_b_75));
SDFFNSRN u9_mem_reg_b3_b_b21_b (.CK(clk_i), .D(n_10710), .Q(u9_mem_b3_b_77), .SO(u9_mem_b3_b_77), .SE(scan_enable), .SI(u9_mem_b3_b_76));
SDFFNSRN u9_mem_reg_b3_b_b23_b (.CK(clk_i), .D(n_10708), .Q(u9_mem_b3_b_79), .SO(u9_mem_b3_b_79), .SE(scan_enable), .SI(u9_mem_b3_b_77));
SDFFNSRN u9_mem_reg_b3_b_b24_b (.CK(clk_i), .D(n_10707), .Q(u9_mem_b3_b_80), .SO(u9_mem_b3_b_80), .SE(scan_enable), .SI(u9_mem_b3_b_79));
SDFFNSRN u9_mem_reg_b3_b_b25_b (.CK(clk_i), .D(n_10706), .Q(u9_mem_b3_b_81), .SO(u9_mem_b3_b_81), .SE(scan_enable), .SI(u9_mem_b3_b_80));
SDFFNSRN u9_mem_reg_b3_b_b27_b (.CK(clk_i), .D(n_10704), .Q(u9_mem_b3_b_83), .SO(u9_mem_b3_b_83), .SE(scan_enable), .SI(u9_mem_b3_b_81));
SDFFNSRN u9_mem_reg_b3_b_b28_b (.CK(clk_i), .D(n_10703), .Q(u9_mem_b3_b_84), .SO(u9_mem_b3_b_84), .SE(scan_enable), .SI(u9_mem_b3_b_83));
SDFFNSRN u9_mem_reg_b3_b_b29_b (.CK(clk_i), .D(n_10702), .Q(u9_mem_b3_b_85), .SO(u9_mem_b3_b_85), .SE(scan_enable), .SI(u9_mem_b3_b_84));
SDFFNSRN u9_mem_reg_b3_b_b31_b (.CK(clk_i), .D(n_10700), .Q(u9_mem_b3_b_87), .SO(u9_mem_b3_b_87), .SE(scan_enable), .SI(u9_mem_b3_b_85));
SDFFNSRN u10_mem_reg_b3_b_b18_b (.CK(clk_i), .D(n_10699), .Q(u10_mem_b3_b_74), .SO(u10_mem_b3_b_74), .SE(scan_enable), .SI(u9_mem_b3_b_87));
SDFFNSRN u10_mem_reg_b3_b_b19_b (.CK(clk_i), .D(n_10697), .Q(u10_mem_b3_b_75), .SO(u10_mem_b3_b_75), .SE(scan_enable), .SI(u10_mem_b3_b_74));
SDFFNSRN u10_mem_reg_b3_b_b20_b (.CK(clk_i), .D(n_10695), .Q(u10_mem_b3_b_76), .SO(u10_mem_b3_b_76), .SE(scan_enable), .SI(u10_mem_b3_b_75));
SDFFNSRN u10_mem_reg_b3_b_b21_b (.CK(clk_i), .D(n_10694), .Q(u10_mem_b3_b_77), .SO(u10_mem_b3_b_77), .SE(scan_enable), .SI(u10_mem_b3_b_76));
SDFFNSRN u10_mem_reg_b3_b_b22_b (.CK(clk_i), .D(n_10693), .Q(u10_mem_b3_b_78), .SO(u10_mem_b3_b_78), .SE(scan_enable), .SI(u10_mem_b3_b_77));
SDFFNSRN u10_mem_reg_b3_b_b23_b (.CK(clk_i), .D(n_10691), .Q(u10_mem_b3_b_79), .SO(u10_mem_b3_b_79), .SE(scan_enable), .SI(u10_mem_b3_b_78));
SDFFNSRN u10_mem_reg_b3_b_b25_b (.CK(clk_i), .D(n_10688), .Q(u10_mem_b3_b_81), .SO(u10_mem_b3_b_81), .SE(scan_enable), .SI(u10_mem_b3_b_79));
SDFFNSRN u10_mem_reg_b3_b_b26_b (.CK(clk_i), .D(n_10686), .Q(u10_mem_b3_b_82), .SO(u10_mem_b3_b_82), .SE(scan_enable), .SI(u10_mem_b3_b_81));
SDFFNSRN u10_mem_reg_b3_b_b27_b (.CK(clk_i), .D(n_10685), .Q(u10_mem_b3_b_83), .SO(u10_mem_b3_b_83), .SE(scan_enable), .SI(u10_mem_b3_b_82));
SDFFNSRN u10_mem_reg_b3_b_b29_b (.CK(clk_i), .D(n_10682), .Q(u10_mem_b3_b_85), .SO(u10_mem_b3_b_85), .SE(scan_enable), .SI(u10_mem_b3_b_83));
SDFFNSRN u10_mem_reg_b3_b_b30_b (.CK(clk_i), .D(n_10681), .Q(u10_mem_b3_b_86), .SO(u10_mem_b3_b_86), .SE(scan_enable), .SI(u10_mem_b3_b_85));
SDFFNSRN u10_mem_reg_b3_b_b31_b (.CK(clk_i), .D(n_10680), .Q(u10_mem_b3_b_87), .SO(u10_mem_b3_b_87), .SE(scan_enable), .SI(u10_mem_b3_b_86));
SDFFNSRN u10_mem_reg_b0_b_b19_b (.CK(clk_i), .D(n_10677), .Q(u10_mem_b0_b_168), .SO(u10_mem_b0_b_168), .SE(scan_enable), .SI(u10_mem_b3_b_87));
SDFFNSRN u10_mem_reg_b1_b_b18_b (.CK(clk_i), .D(n_10676), .Q(u10_mem_b1_b_136), .SO(u10_mem_b1_b_136), .SE(scan_enable), .SI(u10_mem_b0_b_168));
SDFFNSRN u10_mem_reg_b1_b_b19_b (.CK(clk_i), .D(n_10675), .Q(u10_mem_b1_b_137), .SO(u10_mem_b1_b_137), .SE(scan_enable), .SI(u10_mem_b1_b_136));
SDFFNSRN u10_mem_reg_b1_b_b21_b (.CK(clk_i), .D(n_10673), .Q(u10_mem_b1_b_139), .SO(u10_mem_b1_b_139), .SE(scan_enable), .SI(u10_mem_b1_b_137));
SDFFNSRN u10_mem_reg_b1_b_b22_b (.CK(clk_i), .D(n_10672), .Q(u10_mem_b1_b_140), .SO(u10_mem_b1_b_140), .SE(scan_enable), .SI(u10_mem_b1_b_139));
SDFFNSRN u10_mem_reg_b1_b_b23_b (.CK(clk_i), .D(n_10671), .Q(u10_mem_b1_b_141), .SO(u10_mem_b1_b_141), .SE(scan_enable), .SI(u10_mem_b1_b_140));
SDFFNSRN u10_mem_reg_b1_b_b24_b (.CK(clk_i), .D(n_10670), .Q(u10_mem_b1_b_142), .SO(u10_mem_b1_b_142), .SE(scan_enable), .SI(u10_mem_b1_b_141));
SDFFNSRN u10_mem_reg_b1_b_b25_b (.CK(clk_i), .D(n_10669), .Q(u10_mem_b1_b_143), .SO(u10_mem_b1_b_143), .SE(scan_enable), .SI(u10_mem_b1_b_142));
SDFFNSRN u10_mem_reg_b1_b_b26_b (.CK(clk_i), .D(n_10805), .Q(u10_mem_b1_b_144), .SO(u10_mem_b1_b_144), .SE(scan_enable), .SI(u10_mem_b1_b_143));
SDFFNSRN u10_mem_reg_b1_b_b27_b (.CK(clk_i), .D(n_10667), .Q(u10_mem_b1_b_145), .SO(u10_mem_b1_b_145), .SE(scan_enable), .SI(u10_mem_b1_b_144));
SDFFNSRN u10_mem_reg_b1_b_b28_b (.CK(clk_i), .D(n_10666), .Q(u10_mem_b1_b_146), .SO(u10_mem_b1_b_146), .SE(scan_enable), .SI(u10_mem_b1_b_145));
SDFFNSRN u10_mem_reg_b1_b_b29_b (.CK(clk_i), .D(n_10668), .Q(u10_mem_b1_b_147), .SO(u10_mem_b1_b_147), .SE(scan_enable), .SI(u10_mem_b1_b_146));
SDFFNSRN u10_mem_reg_b1_b_b20_b (.CK(clk_i), .D(n_10674), .Q(u10_mem_b1_b_138), .SO(u10_mem_b1_b_138), .SE(scan_enable), .SI(u10_mem_b1_b_147));
SDFFNSRN u10_mem_reg_b1_b_b30_b (.CK(clk_i), .D(n_10664), .Q(u10_mem_b1_b_148), .SO(u10_mem_b1_b_148), .SE(scan_enable), .SI(u10_mem_b1_b_138));
SDFFNSRN u10_mem_reg_b1_b_b31_b (.CK(clk_i), .D(n_10665), .Q(u10_mem_b1_b_149), .SO(u10_mem_b1_b_149), .SE(scan_enable), .SI(u10_mem_b1_b_148));
SDFFNSRN u11_mem_reg_b3_b_b8_b (.CK(clk_i), .D(n_10655), .Q(u11_mem_b3_b_64), .SO(u11_mem_b3_b_64), .SE(scan_enable), .SI(u10_mem_b1_b_149));
SDFFNSRN u11_mem_reg_b3_b_b9_b (.CK(clk_i), .D(n_10654), .Q(u11_mem_b3_b_65), .SO(u11_mem_b3_b_65), .SE(scan_enable), .SI(u11_mem_b3_b_64));
SDFFNSRN u10_mem_reg_b2_b_b1_b (.CK(clk_i), .D(n_10652), .Q(u10_mem_b2_b_88), .SO(u10_mem_b2_b_88), .SE(scan_enable), .SI(u11_mem_b3_b_65));
SDFFNSRN u10_mem_reg_b2_b_b5_b (.CK(clk_i), .D(n_10651), .Q(u10_mem_b2_b_92), .SO(u10_mem_b2_b_92), .SE(scan_enable), .SI(u10_mem_b2_b_88));
SDFFNSRN u10_mem_reg_b2_b_b6_b (.CK(clk_i), .D(n_10649), .Q(u10_mem_b2_b_93), .SO(u10_mem_b2_b_93), .SE(scan_enable), .SI(u10_mem_b2_b_92));
SDFFNSRN u10_mem_reg_b3_b_b3_b (.CK(clk_i), .D(n_10566), .Q(u10_mem_b3_b_59), .SO(u10_mem_b3_b_59), .SE(scan_enable), .SI(u10_mem_b2_b_93));
SDFFNSRN u10_mem_reg_b2_b_b9_b (.CK(clk_i), .D(n_10600), .Q(u10_mem_b2_b_96), .SO(u10_mem_b2_b_96), .SE(scan_enable), .SI(u10_mem_b3_b_59));
SDFFNSRN u11_mem_reg_b1_b_b0_b (.CK(clk_i), .D(n_10563), .Q(u11_mem_b1_b), .SO(u11_mem_b1_b), .SE(scan_enable), .SI(u10_mem_b2_b_96));
SDFFNSRN u11_mem_reg_b1_b_b10_b (.CK(clk_i), .D(n_10562), .Q(u11_mem_b1_b_128), .SO(u11_mem_b1_b_128), .SE(scan_enable), .SI(u11_mem_b1_b));
SDFFNSRN u11_mem_reg_b1_b_b11_b (.CK(clk_i), .D(n_10561), .Q(u11_mem_b1_b_129), .SO(u11_mem_b1_b_129), .SE(scan_enable), .SI(u11_mem_b1_b_128));
SDFFNSRN u10_mem_reg_b3_b_b2_b (.CK(clk_i), .D(n_10567), .Q(u10_mem_b3_b_58), .SO(u10_mem_b3_b_58), .SE(scan_enable), .SI(u11_mem_b1_b_129));
SDFFNSRN u10_mem_reg_b3_b_b9_b (.CK(clk_i), .D(n_10564), .Q(u10_mem_b3_b_65), .SO(u10_mem_b3_b_65), .SE(scan_enable), .SI(u10_mem_b3_b_58));
SDFFNSRN u11_mem_reg_b1_b_b14_b (.CK(clk_i), .D(n_10559), .Q(u11_mem_b1_b_132), .SO(u11_mem_b1_b_132), .SE(scan_enable), .SI(u10_mem_b3_b_65));
SDFFNSRN u11_mem_reg_b1_b_b1_b (.CK(clk_i), .D(n_10555), .Q(u11_mem_b1_b_119), .SO(u11_mem_b1_b_119), .SE(scan_enable), .SI(u11_mem_b1_b_132));
SDFFNSRN u11_mem_reg_b1_b_b2_b (.CK(clk_i), .D(n_10554), .Q(u11_mem_b1_b_120), .SO(u11_mem_b1_b_120), .SE(scan_enable), .SI(u11_mem_b1_b_119));
SDFFNSRN u11_mem_reg_b1_b_b3_b (.CK(clk_i), .D(n_10552), .Q(u11_mem_b1_b_121), .SO(u11_mem_b1_b_121), .SE(scan_enable), .SI(u11_mem_b1_b_120));
SDFFNSRN u11_mem_reg_b1_b_b4_b (.CK(clk_i), .D(n_10551), .Q(u11_mem_b1_b_122), .SO(u11_mem_b1_b_122), .SE(scan_enable), .SI(u11_mem_b1_b_121));
SDFFNSRN u11_mem_reg_b1_b_b5_b (.CK(clk_i), .D(n_10549), .Q(u11_mem_b1_b_123), .SO(u11_mem_b1_b_123), .SE(scan_enable), .SI(u11_mem_b1_b_122));
SDFFNSRN u11_mem_reg_b1_b_b7_b (.CK(clk_i), .D(n_10546), .Q(u11_mem_b1_b_125), .SO(u11_mem_b1_b_125), .SE(scan_enable), .SI(u11_mem_b1_b_123));
SDFFNSRN u11_mem_reg_b1_b_b8_b (.CK(clk_i), .D(n_10545), .Q(u11_mem_b1_b_126), .SO(u11_mem_b1_b_126), .SE(scan_enable), .SI(u11_mem_b1_b_125));
SDFFNSRN u11_mem_reg_b1_b_b9_b (.CK(clk_i), .D(n_10543), .Q(u11_mem_b1_b_127), .SO(u11_mem_b1_b_127), .SE(scan_enable), .SI(u11_mem_b1_b_126));
SDFFNSRN u11_mem_reg_b2_b_b0_b (.CK(clk_i), .D(n_10542), .Q(u11_mem_b2_b), .SO(u11_mem_b2_b), .SE(scan_enable), .SI(u11_mem_b1_b_127));
SDFFNSRN u11_mem_reg_b2_b_b10_b (.CK(clk_i), .D(n_10540), .Q(u11_mem_b2_b_97), .SO(u11_mem_b2_b_97), .SE(scan_enable), .SI(u11_mem_b2_b));
SDFFNSRN u11_mem_reg_b2_b_b11_b (.CK(clk_i), .D(n_10539), .Q(u11_mem_b2_b_98), .SO(u11_mem_b2_b_98), .SE(scan_enable), .SI(u11_mem_b2_b_97));
SDFFNSRN u11_mem_reg_b2_b_b13_b (.CK(clk_i), .D(n_10535), .Q(u11_mem_b2_b_100), .SO(u11_mem_b2_b_100), .SE(scan_enable), .SI(u11_mem_b2_b_98));
SDFFNSRN u11_mem_reg_b2_b_b14_b (.CK(clk_i), .D(n_10529), .Q(u11_mem_b2_b_101), .SO(u11_mem_b2_b_101), .SE(scan_enable), .SI(u11_mem_b2_b_100));
SDFFNSRN u11_mem_reg_b2_b_b15_b (.CK(clk_i), .D(n_10521), .Q(u11_mem_b2_b_102), .SO(u11_mem_b2_b_102), .SE(scan_enable), .SI(u11_mem_b2_b_101));
SDFFNSRN u11_mem_reg_b2_b_b16_b (.CK(clk_i), .D(n_10514), .Q(u11_mem_b2_b_103), .SO(u11_mem_b2_b_103), .SE(scan_enable), .SI(u11_mem_b2_b_102));
SDFFNSRN u11_mem_reg_b1_b_b17_b (.CK(clk_i), .D(n_10556), .Q(u11_mem_b1_b_135), .SO(u11_mem_b1_b_135), .SE(scan_enable), .SI(u11_mem_b2_b_103));
SDFFNSRN u11_mem_reg_b2_b_b12_b (.CK(clk_i), .D(n_10538), .Q(u11_mem_b2_b_99), .SO(u11_mem_b2_b_99), .SE(scan_enable), .SI(u11_mem_b1_b_135));
SDFFNSRN u11_mem_reg_b2_b_b2_b (.CK(clk_i), .D(n_10508), .Q(u11_mem_b2_b_89), .SO(u11_mem_b2_b_89), .SE(scan_enable), .SI(u11_mem_b2_b_99));
SDFFNSRN u11_mem_reg_b2_b_b3_b (.CK(clk_i), .D(n_10501), .Q(u11_mem_b2_b_90), .SO(u11_mem_b2_b_90), .SE(scan_enable), .SI(u11_mem_b2_b_89));
SDFFNSRN u11_mem_reg_b2_b_b6_b (.CK(clk_i), .D(n_10489), .Q(u11_mem_b2_b_93), .SO(u11_mem_b2_b_93), .SE(scan_enable), .SI(u11_mem_b2_b_90));
SDFFNSRN u11_mem_reg_b2_b_b4_b (.CK(clk_i), .D(n_10498), .Q(u11_mem_b2_b_91), .SO(u11_mem_b2_b_91), .SE(scan_enable), .SI(u11_mem_b2_b_93));
SDFFNSRN u11_mem_reg_b2_b_b5_b (.CK(clk_i), .D(n_10494), .Q(u11_mem_b2_b_92), .SO(u11_mem_b2_b_92), .SE(scan_enable), .SI(u11_mem_b2_b_91));
SDFFNSRN u11_mem_reg_b2_b_b9_b (.CK(clk_i), .D(n_10476), .Q(u11_mem_b2_b_96), .SO(u11_mem_b2_b_96), .SE(scan_enable), .SI(u11_mem_b2_b_92));
SDFFNSRN u11_mem_reg_b3_b_b11_b (.CK(clk_i), .D(n_10462), .Q(u11_mem_b3_b_67), .SO(u11_mem_b3_b_67), .SE(scan_enable), .SI(u11_mem_b2_b_96));
SDFFNSRN u11_mem_reg_b3_b_b12_b (.CK(clk_i), .D(n_10459), .Q(u11_mem_b3_b_68), .SO(u11_mem_b3_b_68), .SE(scan_enable), .SI(u11_mem_b3_b_67));
SDFFNSRN u11_mem_reg_b3_b_b15_b (.CK(clk_i), .D(n_10456), .Q(u11_mem_b3_b_71), .SO(u11_mem_b3_b_71), .SE(scan_enable), .SI(u11_mem_b3_b_68));
SDFFNSRN u11_mem_reg_b3_b_b10_b (.CK(clk_i), .D(n_10466), .Q(u11_mem_b3_b_66), .SO(u11_mem_b3_b_66), .SE(scan_enable), .SI(u11_mem_b3_b_71));
SDFFNSRN u11_mem_reg_b3_b_b2_b (.CK(clk_i), .D(n_10454), .Q(u11_mem_b3_b_58), .SO(u11_mem_b3_b_58), .SE(scan_enable), .SI(u11_mem_b3_b_66));
SDFFNSRN u11_mem_reg_b3_b_b3_b (.CK(clk_i), .D(n_10453), .Q(u11_mem_b3_b_59), .SO(u11_mem_b3_b_59), .SE(scan_enable), .SI(u11_mem_b3_b_58));
SDFFNSRN u11_mem_reg_b3_b_b4_b (.CK(clk_i), .D(n_10452), .Q(u11_mem_b3_b_60), .SO(u11_mem_b3_b_60), .SE(scan_enable), .SI(u11_mem_b3_b_59));
SDFFNSRN u11_mem_reg_b3_b_b1_b (.CK(clk_i), .D(n_10455), .Q(u11_mem_b3_b_57), .SO(u11_mem_b3_b_57), .SE(scan_enable), .SI(u11_mem_b3_b_60));
SDFFNSRN u10_wp_reg_b1_b (.CK(clk_i), .D(n_10780), .Q(u10_wp_b1_b), .SO(u10_wp_b1_b), .SE(scan_enable), .SI(u11_mem_b3_b_57));
SDFFNSRN u10_wp_reg_b2_b (.CK(clk_i), .D(n_10801), .Q(u10_wp_b2_b), .SO(u10_wp_b2_b), .SE(scan_enable), .SI(u10_wp_b1_b));
SDFFNSRN u10_mem_reg_b0_b_b2_b (.CK(clk_i), .D(n_10412), .Q(u10_mem_b0_b_151), .SO(u10_mem_b0_b_151), .SE(scan_enable), .SI(u10_wp_b2_b));
SDFFNSRN u11_mem_reg_b0_b_b5_b (.CK(clk_i), .D(n_10422), .Q(u11_mem_b0_b_154), .SO(u11_mem_b0_b_154), .SE(scan_enable), .SI(u10_mem_b0_b_151));
SDFFNSRN u10_mem_reg_b0_b_b13_b (.CK(clk_i), .D(n_10449), .Q(u10_mem_b0_b_162), .SO(u10_mem_b0_b_162), .SE(scan_enable), .SI(u11_mem_b0_b_154));
SDFFNSRN u10_mem_reg_b0_b_b12_b (.CK(clk_i), .D(n_10451), .Q(u10_mem_b0_b_161), .SO(u10_mem_b0_b_161), .SE(scan_enable), .SI(u10_mem_b0_b_162));
SDFFNSRN u11_mem_reg_b0_b_b16_b (.CK(clk_i), .D(n_10448), .Q(u11_mem_b0_b_165), .SO(u11_mem_b0_b_165), .SE(scan_enable), .SI(u10_mem_b0_b_161));
SDFFNSRN u11_mem_reg_b0_b_b20_b (.CK(clk_i), .D(n_10445), .Q(u11_mem_b0_b_169), .SO(u11_mem_b0_b_169), .SE(scan_enable), .SI(u11_mem_b0_b_165));
SDFFNSRN u11_mem_reg_b0_b_b21_b (.CK(clk_i), .D(n_10444), .Q(u11_mem_b0_b_170), .SO(u11_mem_b0_b_170), .SE(scan_enable), .SI(u11_mem_b0_b_169));
SDFFNSRN u11_mem_reg_b0_b_b22_b (.CK(clk_i), .D(n_10443), .Q(u11_mem_b0_b_171), .SO(u11_mem_b0_b_171), .SE(scan_enable), .SI(u11_mem_b0_b_170));
SDFFNSRN u11_mem_reg_b0_b_b23_b (.CK(clk_i), .D(n_10441), .Q(u11_mem_b0_b_172), .SO(u11_mem_b0_b_172), .SE(scan_enable), .SI(u11_mem_b0_b_171));
SDFFNSRN u11_mem_reg_b0_b_b24_b (.CK(clk_i), .D(n_10440), .Q(u11_mem_b0_b_173), .SO(u11_mem_b0_b_173), .SE(scan_enable), .SI(u11_mem_b0_b_172));
SDFFNSRN u11_mem_reg_b0_b_b25_b (.CK(clk_i), .D(n_10439), .Q(u11_mem_b0_b_174), .SO(u11_mem_b0_b_174), .SE(scan_enable), .SI(u11_mem_b0_b_173));
SDFFNSRN u10_mem_reg_b0_b_b21_b (.CK(clk_i), .D(n_10438), .Q(u10_mem_b0_b_170), .SO(u10_mem_b0_b_170), .SE(scan_enable), .SI(u11_mem_b0_b_174));
SDFFNSRN u11_mem_reg_b0_b_b26_b (.CK(clk_i), .D(n_10437), .Q(u11_mem_b0_b_175), .SO(u11_mem_b0_b_175), .SE(scan_enable), .SI(u10_mem_b0_b_170));
SDFFNSRN u11_mem_reg_b0_b_b27_b (.CK(clk_i), .D(n_10436), .Q(u11_mem_b0_b_176), .SO(u11_mem_b0_b_176), .SE(scan_enable), .SI(u11_mem_b0_b_175));
SDFFNSRN u10_mem_reg_b0_b_b22_b (.CK(clk_i), .D(n_10435), .Q(u10_mem_b0_b_171), .SO(u10_mem_b0_b_171), .SE(scan_enable), .SI(u11_mem_b0_b_176));
SDFFNSRN u11_mem_reg_b0_b_b28_b (.CK(clk_i), .D(n_10433), .Q(u11_mem_b0_b_177), .SO(u11_mem_b0_b_177), .SE(scan_enable), .SI(u10_mem_b0_b_171));
SDFFNSRN u11_mem_reg_b0_b_b29_b (.CK(clk_i), .D(n_10432), .Q(u11_mem_b0_b_178), .SO(u11_mem_b0_b_178), .SE(scan_enable), .SI(u11_mem_b0_b_177));
SDFFNSRN u11_mem_reg_b0_b_b2_b (.CK(clk_i), .D(n_10430), .Q(u11_mem_b0_b_151), .SO(u11_mem_b0_b_151), .SE(scan_enable), .SI(u11_mem_b0_b_178));
SDFFNSRN u11_mem_reg_b0_b_b30_b (.CK(clk_i), .D(n_10429), .Q(u11_mem_b0_b_179), .SO(u11_mem_b0_b_179), .SE(scan_enable), .SI(u11_mem_b0_b_151));
SDFFNSRN u11_mem_reg_b0_b_b31_b (.CK(clk_i), .D(n_10428), .Q(u11_mem_b0_b_180), .SO(u11_mem_b0_b_180), .SE(scan_enable), .SI(u11_mem_b0_b_179));
SDFFNSRN u11_mem_reg_b0_b_b3_b (.CK(clk_i), .D(n_10425), .Q(u11_mem_b0_b_152), .SO(u11_mem_b0_b_152), .SE(scan_enable), .SI(u11_mem_b0_b_180));
SDFFNSRN u10_mem_reg_b0_b_b25_b (.CK(clk_i), .D(n_10426), .Q(u10_mem_b0_b_174), .SO(u10_mem_b0_b_174), .SE(scan_enable), .SI(u11_mem_b0_b_152));
SDFFNSRN u11_mem_reg_b0_b_b4_b (.CK(clk_i), .D(n_10424), .Q(u11_mem_b0_b_153), .SO(u11_mem_b0_b_153), .SE(scan_enable), .SI(u10_mem_b0_b_174));
SDFFNSRN u10_mem_reg_b0_b_b26_b (.CK(clk_i), .D(n_10423), .Q(u10_mem_b0_b_175), .SO(u10_mem_b0_b_175), .SE(scan_enable), .SI(u11_mem_b0_b_153));
SDFFNSRN u10_mem_reg_b0_b_b27_b (.CK(clk_i), .D(n_10421), .Q(u10_mem_b0_b_176), .SO(u10_mem_b0_b_176), .SE(scan_enable), .SI(u10_mem_b0_b_175));
SDFFNSRN u11_mem_reg_b0_b_b6_b (.CK(clk_i), .D(n_10420), .Q(u11_mem_b0_b_155), .SO(u11_mem_b0_b_155), .SE(scan_enable), .SI(u10_mem_b0_b_176));
SDFFNSRN u10_mem_reg_b0_b_b28_b (.CK(clk_i), .D(n_10418), .Q(u10_mem_b0_b_177), .SO(u10_mem_b0_b_177), .SE(scan_enable), .SI(u11_mem_b0_b_155));
SDFFNSRN u11_mem_reg_b0_b_b7_b (.CK(clk_i), .D(n_10417), .Q(u11_mem_b0_b_156), .SO(u11_mem_b0_b_156), .SE(scan_enable), .SI(u10_mem_b0_b_177));
SDFFNSRN u11_mem_reg_b0_b_b8_b (.CK(clk_i), .D(n_10416), .Q(u11_mem_b0_b_157), .SO(u11_mem_b0_b_157), .SE(scan_enable), .SI(u11_mem_b0_b_156));
SDFFNSRN u10_mem_reg_b0_b_b29_b (.CK(clk_i), .D(n_10415), .Q(u10_mem_b0_b_178), .SO(u10_mem_b0_b_178), .SE(scan_enable), .SI(u11_mem_b0_b_157));
SDFFNSRN u11_mem_reg_b0_b_b9_b (.CK(clk_i), .D(n_10413), .Q(u11_mem_b0_b_158), .SO(u11_mem_b0_b_158), .SE(scan_enable), .SI(u10_mem_b0_b_178));
SDFFNSRN u10_mem_reg_b0_b_b5_b (.CK(clk_i), .D(n_10411), .Q(u10_mem_b0_b_154), .SO(u10_mem_b0_b_154), .SE(scan_enable), .SI(u11_mem_b0_b_158));
SDFFN u11_wp_reg_b0_b (.CK(clk_i), .D(n_10777), .Q(u11_wp_b0_b), .SO(u11_wp_b0_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u10_mem_b0_b_154));
SDFFN u25_int_set_reg_b2_b (.CK(clk_i), .D(n_10794), .Q(ic2_int_set_724), .SO(ic2_int_set_724), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u11_wp_b0_b));
SDFFNSRN u10_mem_reg_b0_b_b1_b (.CK(clk_i), .D(n_10446), .Q(u10_mem_b0_b_150), .SO(u10_mem_b0_b_150), .SE(scan_enable), .SI(ic2_int_set_724));
SDFFNSRN u11_mem_reg_b0_b_b17_b (.CK(clk_i), .D(n_10447), .Q(u11_mem_b0_b_166), .SO(u11_mem_b0_b_166), .SE(scan_enable), .SI(u10_mem_b0_b_150));
SDFFNSRN u10_mem_reg_b3_b_b17_b (.CK(clk_i), .D(n_10224), .Q(u10_mem_b3_b_73), .SO(u10_mem_b3_b_73), .SE(scan_enable), .SI(u11_mem_b0_b_166));
SDFFNSRN u10_mem_reg_b0_b_b11_b (.CK(clk_i), .D(n_10135), .Q(u10_mem_b0_b_160), .SO(u10_mem_b0_b_160), .SE(scan_enable), .SI(u10_mem_b3_b_73));
SDFFNSRN u9_mem_reg_b0_b_b4_b (.CK(clk_i), .D(n_10147), .Q(u9_mem_b0_b_153), .SO(u9_mem_b0_b_153), .SE(scan_enable), .SI(u10_mem_b0_b_160));
SDFFNSRN u9_wp_reg_b3_b (.CK(clk_i), .D(n_10335), .Q(u9_wp_b3_b), .SO(u9_wp_b3_b), .SE(scan_enable), .SI(u9_mem_b0_b_153));
SDFFNSRN u9_mem_reg_b0_b_b8_b (.CK(clk_i), .D(n_10142), .Q(u9_mem_b0_b_157), .SO(u9_mem_b0_b_157), .SE(scan_enable), .SI(u9_wp_b3_b));
SDFFNSRN u10_mem_reg_b1_b_b8_b (.CK(clk_i), .D(n_10179), .Q(u10_mem_b1_b_126), .SO(u10_mem_b1_b_126), .SE(scan_enable), .SI(u9_mem_b0_b_157));
SDFFNSRN u9_mem_reg_b0_b_b2_b (.CK(clk_i), .D(n_10152), .Q(u9_mem_b0_b_151), .SO(u9_mem_b0_b_151), .SE(scan_enable), .SI(u10_mem_b1_b_126));
SDFFNSRN u9_mem_reg_b0_b_b26_b (.CK(clk_i), .D(n_10157), .Q(u9_mem_b0_b_175), .SO(u9_mem_b0_b_175), .SE(scan_enable), .SI(u9_mem_b0_b_151));
SDFFNSRN u10_mem_reg_b1_b_b6_b (.CK(clk_i), .D(n_10181), .Q(u10_mem_b1_b_124), .SO(u10_mem_b1_b_124), .SE(scan_enable), .SI(u9_mem_b0_b_175));
SDFFNSRN u9_mem_reg_b0_b_b17_b (.CK(clk_i), .D(n_10166), .Q(u9_mem_b0_b_166), .SO(u9_mem_b0_b_166), .SE(scan_enable), .SI(u10_mem_b1_b_124));
SDFFNSRN u9_mem_reg_b0_b_b13_b (.CK(clk_i), .D(n_10170), .Q(u9_mem_b0_b_162), .SO(u9_mem_b0_b_162), .SE(scan_enable), .SI(u9_mem_b0_b_166));
SDFFNSRN u10_mem_reg_b1_b_b1_b (.CK(clk_i), .D(n_10187), .Q(u10_mem_b1_b_119), .SO(u10_mem_b1_b_119), .SE(scan_enable), .SI(u9_mem_b0_b_162));
SDFFNSRN u10_mem_reg_b1_b_b15_b (.CK(clk_i), .D(n_10197), .Q(u10_mem_b1_b_133), .SO(u10_mem_b1_b_133), .SE(scan_enable), .SI(u10_mem_b1_b_119));
SDFFNSRN u10_mem_reg_b1_b_b13_b (.CK(clk_i), .D(n_10211), .Q(u10_mem_b1_b_131), .SO(u10_mem_b1_b_131), .SE(scan_enable), .SI(u10_mem_b1_b_133));
SDFFNSRN u10_mem_reg_b1_b_b10_b (.CK(clk_i), .D(n_10215), .Q(u10_mem_b1_b_128), .SO(u10_mem_b1_b_128), .SE(scan_enable), .SI(u10_mem_b1_b_131));
SDFFNSRN u10_mem_reg_b3_b_b8_b (.CK(clk_i), .D(n_10216), .Q(u10_mem_b3_b_64), .SO(u10_mem_b3_b_64), .SE(scan_enable), .SI(u10_mem_b1_b_128));
SDFFNSRN u10_mem_reg_b0_b_b23_b (.CK(clk_i), .D(n_10129), .Q(u10_mem_b0_b_172), .SO(u10_mem_b0_b_172), .SE(scan_enable), .SI(u10_mem_b3_b_64));
SDFFNSRN u11_din_tmp1_reg_b8_b (.CK(clk_i), .D(n_10097), .Q(u11_din_tmp_49), .SO(u11_din_tmp_49), .SE(scan_enable), .SI(u10_mem_b0_b_172));
SDFFNSRN u9_mem_reg_b2_b_b12_b (.CK(clk_i), .D(n_10285), .Q(u9_mem_b2_b_99), .SO(u9_mem_b2_b_99), .SE(scan_enable), .SI(u11_din_tmp_49));
SDFFNSRN u10_mem_reg_b3_b_b13_b (.CK(clk_i), .D(n_10229), .Q(u10_mem_b3_b_69), .SO(u10_mem_b3_b_69), .SE(scan_enable), .SI(u9_mem_b2_b_99));
SDFFNSRN u10_mem_reg_b3_b_b0_b (.CK(clk_i), .D(n_10234), .Q(u10_mem_b3_b), .SO(u10_mem_b3_b), .SE(scan_enable), .SI(u10_mem_b3_b_69));
SDFFNSRN u9_mem_reg_b3_b_b4_b (.CK(clk_i), .D(n_10243), .Q(u9_mem_b3_b_60), .SO(u9_mem_b3_b_60), .SE(scan_enable), .SI(u10_mem_b3_b));
SDFFNSRN u9_mem_reg_b3_b_b1_b (.CK(clk_i), .D(n_10251), .Q(u9_mem_b3_b_57), .SO(u9_mem_b3_b_57), .SE(scan_enable), .SI(u9_mem_b3_b_60));
SDFFNSRN u9_mem_reg_b3_b_b15_b (.CK(clk_i), .D(n_10254), .Q(u9_mem_b3_b_71), .SO(u9_mem_b3_b_71), .SE(scan_enable), .SI(u9_mem_b3_b_57));
SDFFNSRN u9_mem_reg_b2_b_b5_b (.CK(clk_i), .D(n_10269), .Q(u9_mem_b2_b_92), .SO(u9_mem_b2_b_92), .SE(scan_enable), .SI(u9_mem_b3_b_71));
SDFFNSRN u9_mem_reg_b2_b_b2_b (.CK(clk_i), .D(n_10275), .Q(u9_mem_b2_b_89), .SO(u9_mem_b2_b_89), .SE(scan_enable), .SI(u9_mem_b2_b_92));
SDFFNSRN u10_mem_reg_b1_b_b9_b (.CK(clk_i), .D(n_10178), .Q(u10_mem_b1_b_127), .SO(u10_mem_b1_b_127), .SE(scan_enable), .SI(u9_mem_b2_b_89));
SDFFNSRN u10_mem_reg_b2_b_b0_b (.CK(clk_i), .D(n_10326), .Q(u10_mem_b2_b), .SO(u10_mem_b2_b), .SE(scan_enable), .SI(u10_mem_b1_b_127));
SDFFNSRN u10_mem_reg_b2_b_b11_b (.CK(clk_i), .D(n_10323), .Q(u10_mem_b2_b_98), .SO(u10_mem_b2_b_98), .SE(scan_enable), .SI(u10_mem_b2_b));
SDFFNSRN u10_mem_reg_b2_b_b12_b (.CK(clk_i), .D(n_10322), .Q(u10_mem_b2_b_99), .SO(u10_mem_b2_b_99), .SE(scan_enable), .SI(u10_mem_b2_b_98));
SDFFNSRN u10_mem_reg_b2_b_b13_b (.CK(clk_i), .D(n_10321), .Q(u10_mem_b2_b_100), .SO(u10_mem_b2_b_100), .SE(scan_enable), .SI(u10_mem_b2_b_99));
SDFFNSRN u10_mem_reg_b2_b_b14_b (.CK(clk_i), .D(n_10319), .Q(u10_mem_b2_b_101), .SO(u10_mem_b2_b_101), .SE(scan_enable), .SI(u10_mem_b2_b_100));
SDFFNSRN u10_mem_reg_b2_b_b15_b (.CK(clk_i), .D(n_10318), .Q(u10_mem_b2_b_102), .SO(u10_mem_b2_b_102), .SE(scan_enable), .SI(u10_mem_b2_b_101));
SDFFNSRN u10_mem_reg_b2_b_b16_b (.CK(clk_i), .D(n_10317), .Q(u10_mem_b2_b_103), .SO(u10_mem_b2_b_103), .SE(scan_enable), .SI(u10_mem_b2_b_102));
SDFFNSRN u10_mem_reg_b2_b_b10_b (.CK(clk_i), .D(n_10325), .Q(u10_mem_b2_b_97), .SO(u10_mem_b2_b_97), .SE(scan_enable), .SI(u10_mem_b2_b_103));
SDFFNSRN u9_mem_reg_b1_b_b0_b (.CK(clk_i), .D(n_10314), .Q(u9_mem_b1_b), .SO(u9_mem_b1_b), .SE(scan_enable), .SI(u10_mem_b2_b_97));
SDFFNSRN u9_mem_reg_b1_b_b10_b (.CK(clk_i), .D(n_10313), .Q(u9_mem_b1_b_128), .SO(u9_mem_b1_b_128), .SE(scan_enable), .SI(u9_mem_b1_b));
SDFFNSRN u9_mem_reg_b1_b_b12_b (.CK(clk_i), .D(n_10310), .Q(u9_mem_b1_b_130), .SO(u9_mem_b1_b_130), .SE(scan_enable), .SI(u9_mem_b1_b_128));
SDFFNSRN u9_mem_reg_b1_b_b13_b (.CK(clk_i), .D(n_10309), .Q(u9_mem_b1_b_131), .SO(u9_mem_b1_b_131), .SE(scan_enable), .SI(u9_mem_b1_b_130));
SDFFNSRN u9_mem_reg_b1_b_b14_b (.CK(clk_i), .D(n_10307), .Q(u9_mem_b1_b_132), .SO(u9_mem_b1_b_132), .SE(scan_enable), .SI(u9_mem_b1_b_131));
SDFFNSRN u9_mem_reg_b1_b_b16_b (.CK(clk_i), .D(n_10305), .Q(u9_mem_b1_b_134), .SO(u9_mem_b1_b_134), .SE(scan_enable), .SI(u9_mem_b1_b_132));
SDFFNSRN u9_mem_reg_b1_b_b17_b (.CK(clk_i), .D(n_10304), .Q(u9_mem_b1_b_135), .SO(u9_mem_b1_b_135), .SE(scan_enable), .SI(u9_mem_b1_b_134));
SDFFNSRN u9_mem_reg_b1_b_b1_b (.CK(clk_i), .D(n_10302), .Q(u9_mem_b1_b_119), .SO(u9_mem_b1_b_119), .SE(scan_enable), .SI(u9_mem_b1_b_135));
SDFFNSRN u9_mem_reg_b1_b_b2_b (.CK(clk_i), .D(n_10300), .Q(u9_mem_b1_b_120), .SO(u9_mem_b1_b_120), .SE(scan_enable), .SI(u9_mem_b1_b_119));
SDFFNSRN u9_mem_reg_b1_b_b3_b (.CK(clk_i), .D(n_10299), .Q(u9_mem_b1_b_121), .SO(u9_mem_b1_b_121), .SE(scan_enable), .SI(u9_mem_b1_b_120));
SDFFNSRN u9_mem_reg_b1_b_b4_b (.CK(clk_i), .D(n_10298), .Q(u9_mem_b1_b_122), .SO(u9_mem_b1_b_122), .SE(scan_enable), .SI(u9_mem_b1_b_121));
SDFFNSRN u9_mem_reg_b1_b_b5_b (.CK(clk_i), .D(n_10296), .Q(u9_mem_b1_b_123), .SO(u9_mem_b1_b_123), .SE(scan_enable), .SI(u9_mem_b1_b_122));
SDFFNSRN u9_mem_reg_b1_b_b6_b (.CK(clk_i), .D(n_10295), .Q(u9_mem_b1_b_124), .SO(u9_mem_b1_b_124), .SE(scan_enable), .SI(u9_mem_b1_b_123));
SDFFNSRN u9_mem_reg_b1_b_b7_b (.CK(clk_i), .D(n_10293), .Q(u9_mem_b1_b_125), .SO(u9_mem_b1_b_125), .SE(scan_enable), .SI(u9_mem_b1_b_124));
SDFFNSRN u9_mem_reg_b1_b_b8_b (.CK(clk_i), .D(n_10291), .Q(u9_mem_b1_b_126), .SO(u9_mem_b1_b_126), .SE(scan_enable), .SI(u9_mem_b1_b_125));
SDFFNSRN u9_mem_reg_b2_b_b0_b (.CK(clk_i), .D(n_10289), .Q(u9_mem_b2_b), .SO(u9_mem_b2_b), .SE(scan_enable), .SI(u9_mem_b1_b_126));
SDFFNSRN u9_mem_reg_b2_b_b10_b (.CK(clk_i), .D(n_10288), .Q(u9_mem_b2_b_97), .SO(u9_mem_b2_b_97), .SE(scan_enable), .SI(u9_mem_b2_b));
SDFFNSRN u9_mem_reg_b2_b_b11_b (.CK(clk_i), .D(n_10287), .Q(u9_mem_b2_b_98), .SO(u9_mem_b2_b_98), .SE(scan_enable), .SI(u9_mem_b2_b_97));
SDFFNSRN u9_mem_reg_b2_b_b14_b (.CK(clk_i), .D(n_10283), .Q(u9_mem_b2_b_101), .SO(u9_mem_b2_b_101), .SE(scan_enable), .SI(u9_mem_b2_b_98));
SDFFNSRN u9_mem_reg_b2_b_b15_b (.CK(clk_i), .D(n_10281), .Q(u9_mem_b2_b_102), .SO(u9_mem_b2_b_102), .SE(scan_enable), .SI(u9_mem_b2_b_101));
SDFFNSRN u9_mem_reg_b2_b_b16_b (.CK(clk_i), .D(n_10280), .Q(u9_mem_b2_b_103), .SO(u9_mem_b2_b_103), .SE(scan_enable), .SI(u9_mem_b2_b_102));
SDFFNSRN u9_mem_reg_b2_b_b17_b (.CK(clk_i), .D(n_10279), .Q(u9_mem_b2_b_104), .SO(u9_mem_b2_b_104), .SE(scan_enable), .SI(u9_mem_b2_b_103));
SDFFNSRN u9_mem_reg_b2_b_b1_b (.CK(clk_i), .D(n_10278), .Q(u9_mem_b2_b_88), .SO(u9_mem_b2_b_88), .SE(scan_enable), .SI(u9_mem_b2_b_104));
SDFFNSRN u10_mem_reg_b2_b_b3_b (.CK(clk_i), .D(n_10276), .Q(u10_mem_b2_b_90), .SO(u10_mem_b2_b_90), .SE(scan_enable), .SI(u9_mem_b2_b_88));
SDFFNSRN u9_mem_reg_b2_b_b3_b (.CK(clk_i), .D(n_10272), .Q(u9_mem_b2_b_90), .SO(u9_mem_b2_b_90), .SE(scan_enable), .SI(u10_mem_b2_b_90));
SDFFNSRN u10_mem_reg_b2_b_b4_b (.CK(clk_i), .D(n_10274), .Q(u10_mem_b2_b_91), .SO(u10_mem_b2_b_91), .SE(scan_enable), .SI(u9_mem_b2_b_90));
SDFFNSRN u9_mem_reg_b2_b_b4_b (.CK(clk_i), .D(n_10270), .Q(u9_mem_b2_b_91), .SO(u9_mem_b2_b_91), .SE(scan_enable), .SI(u10_mem_b2_b_91));
SDFFNSRN u9_mem_reg_b2_b_b6_b (.CK(clk_i), .D(n_10268), .Q(u9_mem_b2_b_93), .SO(u9_mem_b2_b_93), .SE(scan_enable), .SI(u9_mem_b2_b_91));
SDFFNSRN u9_mem_reg_b2_b_b7_b (.CK(clk_i), .D(n_10266), .Q(u9_mem_b2_b_94), .SO(u9_mem_b2_b_94), .SE(scan_enable), .SI(u9_mem_b2_b_93));
SDFFNSRN u9_mem_reg_b2_b_b8_b (.CK(clk_i), .D(n_10265), .Q(u9_mem_b2_b_95), .SO(u9_mem_b2_b_95), .SE(scan_enable), .SI(u9_mem_b2_b_94));
SDFFNSRN u9_mem_reg_b3_b_b0_b (.CK(clk_i), .D(n_10263), .Q(u9_mem_b3_b), .SO(u9_mem_b3_b), .SE(scan_enable), .SI(u9_mem_b2_b_95));
SDFFNSRN u9_mem_reg_b3_b_b10_b (.CK(clk_i), .D(n_10262), .Q(u9_mem_b3_b_66), .SO(u9_mem_b3_b_66), .SE(scan_enable), .SI(u9_mem_b3_b));
SDFFNSRN u9_mem_reg_b3_b_b11_b (.CK(clk_i), .D(n_10261), .Q(u9_mem_b3_b_67), .SO(u9_mem_b3_b_67), .SE(scan_enable), .SI(u9_mem_b3_b_66));
SDFFNSRN u9_mem_reg_b3_b_b12_b (.CK(clk_i), .D(n_10259), .Q(u9_mem_b3_b_68), .SO(u9_mem_b3_b_68), .SE(scan_enable), .SI(u9_mem_b3_b_67));
SDFFNSRN u9_mem_reg_b3_b_b13_b (.CK(clk_i), .D(n_10258), .Q(u9_mem_b3_b_69), .SO(u9_mem_b3_b_69), .SE(scan_enable), .SI(u9_mem_b3_b_68));
SDFFNSRN u9_mem_reg_b3_b_b14_b (.CK(clk_i), .D(n_10256), .Q(u9_mem_b3_b_70), .SO(u9_mem_b3_b_70), .SE(scan_enable), .SI(u9_mem_b3_b_69));
SDFFNSRN u9_mem_reg_b2_b_b13_b (.CK(clk_i), .D(n_10284), .Q(u9_mem_b2_b_100), .SO(u9_mem_b2_b_100), .SE(scan_enable), .SI(u9_mem_b3_b_70));
SDFFNSRN u9_mem_reg_b3_b_b16_b (.CK(clk_i), .D(n_10253), .Q(u9_mem_b3_b_72), .SO(u9_mem_b3_b_72), .SE(scan_enable), .SI(u9_mem_b2_b_100));
SDFFNSRN u9_mem_reg_b3_b_b17_b (.CK(clk_i), .D(n_10252), .Q(u9_mem_b3_b_73), .SO(u9_mem_b3_b_73), .SE(scan_enable), .SI(u9_mem_b3_b_72));
SDFFNSRN u10_mem_reg_b2_b_b7_b (.CK(clk_i), .D(n_10249), .Q(u10_mem_b2_b_94), .SO(u10_mem_b2_b_94), .SE(scan_enable), .SI(u9_mem_b3_b_73));
SDFFNSRN u9_mem_reg_b3_b_b2_b (.CK(clk_i), .D(n_10247), .Q(u9_mem_b3_b_58), .SO(u9_mem_b3_b_58), .SE(scan_enable), .SI(u10_mem_b2_b_94));
SDFFNSRN u9_mem_reg_b3_b_b3_b (.CK(clk_i), .D(n_10245), .Q(u9_mem_b3_b_59), .SO(u9_mem_b3_b_59), .SE(scan_enable), .SI(u9_mem_b3_b_58));
SDFFNSRN u9_mem_reg_b3_b_b5_b (.CK(clk_i), .D(n_10242), .Q(u9_mem_b3_b_61), .SO(u9_mem_b3_b_61), .SE(scan_enable), .SI(u9_mem_b3_b_59));
SDFFNSRN u9_mem_reg_b3_b_b6_b (.CK(clk_i), .D(n_10241), .Q(u9_mem_b3_b_62), .SO(u9_mem_b3_b_62), .SE(scan_enable), .SI(u9_mem_b3_b_61));
SDFFNSRN u9_mem_reg_b3_b_b7_b (.CK(clk_i), .D(n_10239), .Q(u9_mem_b3_b_63), .SO(u9_mem_b3_b_63), .SE(scan_enable), .SI(u9_mem_b3_b_62));
SDFFNSRN u10_mem_reg_b2_b_b8_b (.CK(clk_i), .D(n_10244), .Q(u10_mem_b2_b_95), .SO(u10_mem_b2_b_95), .SE(scan_enable), .SI(u9_mem_b3_b_63));
SDFFNSRN u9_mem_reg_b3_b_b9_b (.CK(clk_i), .D(n_10236), .Q(u9_mem_b3_b_65), .SO(u9_mem_b3_b_65), .SE(scan_enable), .SI(u10_mem_b2_b_95));
SDFFNSRN u9_mem_reg_b3_b_b8_b (.CK(clk_i), .D(n_10238), .Q(u9_mem_b3_b_64), .SO(u9_mem_b3_b_64), .SE(scan_enable), .SI(u9_mem_b3_b_65));
SDFFNSRN u10_mem_reg_b3_b_b10_b (.CK(clk_i), .D(n_10233), .Q(u10_mem_b3_b_66), .SO(u10_mem_b3_b_66), .SE(scan_enable), .SI(u9_mem_b3_b_64));
SDFFNSRN u10_mem_reg_b3_b_b11_b (.CK(clk_i), .D(n_10232), .Q(u10_mem_b3_b_67), .SO(u10_mem_b3_b_67), .SE(scan_enable), .SI(u10_mem_b3_b_66));
SDFFNSRN u10_mem_reg_b3_b_b12_b (.CK(clk_i), .D(n_10230), .Q(u10_mem_b3_b_68), .SO(u10_mem_b3_b_68), .SE(scan_enable), .SI(u10_mem_b3_b_67));
SDFFNSRN u10_mem_reg_b3_b_b14_b (.CK(clk_i), .D(n_10228), .Q(u10_mem_b3_b_70), .SO(u10_mem_b3_b_70), .SE(scan_enable), .SI(u10_mem_b3_b_68));
SDFFNSRN u10_mem_reg_b3_b_b15_b (.CK(clk_i), .D(n_10226), .Q(u10_mem_b3_b_71), .SO(u10_mem_b3_b_71), .SE(scan_enable), .SI(u10_mem_b3_b_70));
SDFFNSRN u10_mem_reg_b3_b_b16_b (.CK(clk_i), .D(n_10225), .Q(u10_mem_b3_b_72), .SO(u10_mem_b3_b_72), .SE(scan_enable), .SI(u10_mem_b3_b_71));
SDFFNSRN u10_mem_reg_b3_b_b1_b (.CK(clk_i), .D(n_10223), .Q(u10_mem_b3_b_57), .SO(u10_mem_b3_b_57), .SE(scan_enable), .SI(u10_mem_b3_b_72));
SDFFNSRN u10_mem_reg_b3_b_b4_b (.CK(clk_i), .D(n_10221), .Q(u10_mem_b3_b_60), .SO(u10_mem_b3_b_60), .SE(scan_enable), .SI(u10_mem_b3_b_57));
SDFFNSRN u10_mem_reg_b3_b_b5_b (.CK(clk_i), .D(n_10220), .Q(u10_mem_b3_b_61), .SO(u10_mem_b3_b_61), .SE(scan_enable), .SI(u10_mem_b3_b_60));
SDFFNSRN u10_mem_reg_b3_b_b6_b (.CK(clk_i), .D(n_10219), .Q(u10_mem_b3_b_62), .SO(u10_mem_b3_b_62), .SE(scan_enable), .SI(u10_mem_b3_b_61));
SDFFNSRN u10_mem_reg_b3_b_b7_b (.CK(clk_i), .D(n_10217), .Q(u10_mem_b3_b_63), .SO(u10_mem_b3_b_63), .SE(scan_enable), .SI(u10_mem_b3_b_62));
SDFFNSRN u10_mem_reg_b1_b_b11_b (.CK(clk_i), .D(n_10214), .Q(u10_mem_b1_b_129), .SO(u10_mem_b1_b_129), .SE(scan_enable), .SI(u10_mem_b3_b_63));
SDFFNSRN u10_mem_reg_b1_b_b12_b (.CK(clk_i), .D(n_10212), .Q(u10_mem_b1_b_130), .SO(u10_mem_b1_b_130), .SE(scan_enable), .SI(u10_mem_b1_b_129));
SDFFNSRN u10_mem_reg_b1_b_b14_b (.CK(clk_i), .D(n_10205), .Q(u10_mem_b1_b_132), .SO(u10_mem_b1_b_132), .SE(scan_enable), .SI(u10_mem_b1_b_130));
SDFFNSRN u10_mem_reg_b1_b_b17_b (.CK(clk_i), .D(n_10190), .Q(u10_mem_b1_b_135), .SO(u10_mem_b1_b_135), .SE(scan_enable), .SI(u10_mem_b1_b_132));
SDFFNSRN u10_mem_reg_b1_b_b16_b (.CK(clk_i), .D(n_10194), .Q(u10_mem_b1_b_134), .SO(u10_mem_b1_b_134), .SE(scan_enable), .SI(u10_mem_b1_b_135));
SDFFNSRN u9_mem_reg_b1_b_b9_b (.CK(clk_i), .D(n_10290), .Q(u9_mem_b1_b_127), .SO(u9_mem_b1_b_127), .SE(scan_enable), .SI(u10_mem_b1_b_134));
SDFFNSRN u10_mem_reg_b1_b_b3_b (.CK(clk_i), .D(n_10184), .Q(u10_mem_b1_b_121), .SO(u10_mem_b1_b_121), .SE(scan_enable), .SI(u9_mem_b1_b_127));
SDFFNSRN u10_mem_reg_b1_b_b4_b (.CK(clk_i), .D(n_10183), .Q(u10_mem_b1_b_122), .SO(u10_mem_b1_b_122), .SE(scan_enable), .SI(u10_mem_b1_b_121));
SDFFNSRN u10_mem_reg_b1_b_b5_b (.CK(clk_i), .D(n_10182), .Q(u10_mem_b1_b_123), .SO(u10_mem_b1_b_123), .SE(scan_enable), .SI(u10_mem_b1_b_122));
SDFFNSRN u10_mem_reg_b1_b_b2_b (.CK(clk_i), .D(n_10185), .Q(u10_mem_b1_b_120), .SO(u10_mem_b1_b_120), .SE(scan_enable), .SI(u10_mem_b1_b_123));
SDFFNSRN u10_mem_reg_b2_b_b2_b (.CK(clk_i), .D(n_10301), .Q(u10_mem_b2_b_89), .SO(u10_mem_b2_b_89), .SE(scan_enable), .SI(u10_mem_b1_b_120));
SDFFNSRN u10_mem_reg_b1_b_b7_b (.CK(clk_i), .D(n_10180), .Q(u10_mem_b1_b_125), .SO(u10_mem_b1_b_125), .SE(scan_enable), .SI(u10_mem_b2_b_89));
SDFFNSRN u9_wp_reg_b2_b (.CK(clk_i), .D(n_10394), .Q(u9_wp_b2_b), .SO(u9_wp_b2_b), .SE(scan_enable), .SI(u10_mem_b1_b_125));
SDFFNSRN u9_mem_reg_b1_b_b15_b (.CK(clk_i), .D(n_10306), .Q(u9_mem_b1_b_133), .SO(u9_mem_b1_b_133), .SE(scan_enable), .SI(u9_wp_b2_b));
SDFFNSRN u9_mem_reg_b1_b_b11_b (.CK(clk_i), .D(n_10311), .Q(u9_mem_b1_b_129), .SO(u9_mem_b1_b_129), .SE(scan_enable), .SI(u9_mem_b1_b_133));
SDFFNSRN u10_mem_reg_b2_b_b17_b (.CK(clk_i), .D(n_10316), .Q(u10_mem_b2_b_104), .SO(u10_mem_b2_b_104), .SE(scan_enable), .SI(u9_mem_b1_b_129));
SDFFNSRN u10_mem_reg_b0_b_b24_b (.CK(clk_i), .D(n_10128), .Q(u10_mem_b0_b_173), .SO(u10_mem_b0_b_173), .SE(scan_enable), .SI(u10_mem_b2_b_104));
SDFFNSRN u11_din_tmp1_reg_b4_b (.CK(clk_i), .D(n_10101), .Q(u11_din_tmp_45), .SO(u11_din_tmp_45), .SE(scan_enable), .SI(u10_mem_b0_b_173));
SDFFNSRN u10_mem_reg_b0_b_b8_b (.CK(clk_i), .D(n_10119), .Q(u10_mem_b0_b_157), .SO(u10_mem_b0_b_157), .SE(scan_enable), .SI(u11_din_tmp_45));
SDFFNSRN u10_mem_reg_b0_b_b4_b (.CK(clk_i), .D(n_10123), .Q(u10_mem_b0_b_153), .SO(u10_mem_b0_b_153), .SE(scan_enable), .SI(u10_mem_b0_b_157));
SDFFNSRN u9_mem_reg_b0_b_b0_b (.CK(clk_i), .D(n_10176), .Q(u9_mem_b0_b), .SO(u9_mem_b0_b), .SE(scan_enable), .SI(u10_mem_b0_b_153));
SDFFNSRN u9_mem_reg_b0_b_b10_b (.CK(clk_i), .D(n_10174), .Q(u9_mem_b0_b_159), .SO(u9_mem_b0_b_159), .SE(scan_enable), .SI(u9_mem_b0_b));
SDFFNSRN u9_mem_reg_b0_b_b11_b (.CK(clk_i), .D(n_10173), .Q(u9_mem_b0_b_160), .SO(u9_mem_b0_b_160), .SE(scan_enable), .SI(u9_mem_b0_b_159));
SDFFNSRN u9_mem_reg_b0_b_b12_b (.CK(clk_i), .D(n_10172), .Q(u9_mem_b0_b_161), .SO(u9_mem_b0_b_161), .SE(scan_enable), .SI(u9_mem_b0_b_160));
SDFFNSRN u9_mem_reg_b0_b_b14_b (.CK(clk_i), .D(n_10169), .Q(u9_mem_b0_b_163), .SO(u9_mem_b0_b_163), .SE(scan_enable), .SI(u9_mem_b0_b_161));
SDFFNSRN u9_mem_reg_b0_b_b15_b (.CK(clk_i), .D(n_10168), .Q(u9_mem_b0_b_164), .SO(u9_mem_b0_b_164), .SE(scan_enable), .SI(u9_mem_b0_b_163));
SDFFNSRN u9_mem_reg_b0_b_b16_b (.CK(clk_i), .D(n_10167), .Q(u9_mem_b0_b_165), .SO(u9_mem_b0_b_165), .SE(scan_enable), .SI(u9_mem_b0_b_164));
SDFFNSRN u9_mem_reg_b0_b_b1_b (.CK(clk_i), .D(n_10165), .Q(u9_mem_b0_b_150), .SO(u9_mem_b0_b_150), .SE(scan_enable), .SI(u9_mem_b0_b_165));
SDFFNSRN u9_mem_reg_b0_b_b20_b (.CK(clk_i), .D(n_10164), .Q(u9_mem_b0_b_169), .SO(u9_mem_b0_b_169), .SE(scan_enable), .SI(u9_mem_b0_b_150));
SDFFNSRN u9_mem_reg_b0_b_b21_b (.CK(clk_i), .D(n_10163), .Q(u9_mem_b0_b_170), .SO(u9_mem_b0_b_170), .SE(scan_enable), .SI(u9_mem_b0_b_169));
SDFFNSRN u9_mem_reg_b0_b_b22_b (.CK(clk_i), .D(n_10162), .Q(u9_mem_b0_b_171), .SO(u9_mem_b0_b_171), .SE(scan_enable), .SI(u9_mem_b0_b_170));
SDFFNSRN u9_mem_reg_b0_b_b23_b (.CK(clk_i), .D(n_10160), .Q(u9_mem_b0_b_172), .SO(u9_mem_b0_b_172), .SE(scan_enable), .SI(u9_mem_b0_b_171));
SDFFNSRN u9_mem_reg_b0_b_b24_b (.CK(clk_i), .D(n_10159), .Q(u9_mem_b0_b_173), .SO(u9_mem_b0_b_173), .SE(scan_enable), .SI(u9_mem_b0_b_172));
SDFFNSRN u9_mem_reg_b0_b_b25_b (.CK(clk_i), .D(n_10158), .Q(u9_mem_b0_b_174), .SO(u9_mem_b0_b_174), .SE(scan_enable), .SI(u9_mem_b0_b_173));
SDFFNSRN u9_mem_reg_b0_b_b27_b (.CK(clk_i), .D(n_10156), .Q(u9_mem_b0_b_176), .SO(u9_mem_b0_b_176), .SE(scan_enable), .SI(u9_mem_b0_b_174));
SDFFNSRN u9_mem_reg_b0_b_b28_b (.CK(clk_i), .D(n_10155), .Q(u9_mem_b0_b_177), .SO(u9_mem_b0_b_177), .SE(scan_enable), .SI(u9_mem_b0_b_176));
SDFFNSRN u9_mem_reg_b0_b_b29_b (.CK(clk_i), .D(n_10154), .Q(u9_mem_b0_b_178), .SO(u9_mem_b0_b_178), .SE(scan_enable), .SI(u9_mem_b0_b_177));
SDFFNSRN u9_mem_reg_b0_b_b30_b (.CK(clk_i), .D(n_10151), .Q(u9_mem_b0_b_179), .SO(u9_mem_b0_b_179), .SE(scan_enable), .SI(u9_mem_b0_b_178));
SDFFNSRN u9_mem_reg_b0_b_b31_b (.CK(clk_i), .D(n_10150), .Q(u9_mem_b0_b_180), .SO(u9_mem_b0_b_180), .SE(scan_enable), .SI(u9_mem_b0_b_179));
SDFFNSRN u9_mem_reg_b0_b_b3_b (.CK(clk_i), .D(n_10148), .Q(u9_mem_b0_b_152), .SO(u9_mem_b0_b_152), .SE(scan_enable), .SI(u9_mem_b0_b_180));
SDFFNSRN u9_mem_reg_b0_b_b5_b (.CK(clk_i), .D(n_10146), .Q(u9_mem_b0_b_154), .SO(u9_mem_b0_b_154), .SE(scan_enable), .SI(u9_mem_b0_b_152));
SDFFNSRN u9_mem_reg_b0_b_b6_b (.CK(clk_i), .D(n_10145), .Q(u9_mem_b0_b_155), .SO(u9_mem_b0_b_155), .SE(scan_enable), .SI(u9_mem_b0_b_154));
SDFFNSRN u9_mem_reg_b0_b_b7_b (.CK(clk_i), .D(n_10143), .Q(u9_mem_b0_b_156), .SO(u9_mem_b0_b_156), .SE(scan_enable), .SI(u9_mem_b0_b_155));
SDFFNSRN u9_mem_reg_b0_b_b9_b (.CK(clk_i), .D(n_10141), .Q(u9_mem_b0_b_158), .SO(u9_mem_b0_b_158), .SE(scan_enable), .SI(u9_mem_b0_b_156));
SDFFNSRN u10_mem_reg_b0_b_b0_b (.CK(clk_i), .D(n_10138), .Q(u10_mem_b0_b), .SO(u10_mem_b0_b), .SE(scan_enable), .SI(u9_mem_b0_b_158));
SDFFNSRN u10_mem_reg_b0_b_b10_b (.CK(clk_i), .D(n_10136), .Q(u10_mem_b0_b_159), .SO(u10_mem_b0_b_159), .SE(scan_enable), .SI(u10_mem_b0_b));
SDFFNSRN u10_mem_reg_b0_b_b14_b (.CK(clk_i), .D(n_10134), .Q(u10_mem_b0_b_163), .SO(u10_mem_b0_b_163), .SE(scan_enable), .SI(u10_mem_b0_b_159));
SDFFNSRN u10_mem_reg_b0_b_b15_b (.CK(clk_i), .D(n_10133), .Q(u10_mem_b0_b_164), .SO(u10_mem_b0_b_164), .SE(scan_enable), .SI(u10_mem_b0_b_163));
SDFFNSRN u10_mem_reg_b0_b_b16_b (.CK(clk_i), .D(n_10132), .Q(u10_mem_b0_b_165), .SO(u10_mem_b0_b_165), .SE(scan_enable), .SI(u10_mem_b0_b_164));
SDFFNSRN u10_mem_reg_b0_b_b17_b (.CK(clk_i), .D(n_10131), .Q(u10_mem_b0_b_166), .SO(u10_mem_b0_b_166), .SE(scan_enable), .SI(u10_mem_b0_b_165));
SDFFNSRN u10_mem_reg_b0_b_b31_b (.CK(clk_i), .D(n_10126), .Q(u10_mem_b0_b_180), .SO(u10_mem_b0_b_180), .SE(scan_enable), .SI(u10_mem_b0_b_166));
SDFFNSRN u10_mem_reg_b0_b_b3_b (.CK(clk_i), .D(n_10124), .Q(u10_mem_b0_b_152), .SO(u10_mem_b0_b_152), .SE(scan_enable), .SI(u10_mem_b0_b_180));
SDFFNSRN u10_mem_reg_b0_b_b30_b (.CK(clk_i), .D(n_10127), .Q(u10_mem_b0_b_179), .SO(u10_mem_b0_b_179), .SE(scan_enable), .SI(u10_mem_b0_b_152));
SDFFNSRN u10_mem_reg_b0_b_b6_b (.CK(clk_i), .D(n_10122), .Q(u10_mem_b0_b_155), .SO(u10_mem_b0_b_155), .SE(scan_enable), .SI(u10_mem_b0_b_179));
SDFFNSRN u10_mem_reg_b0_b_b7_b (.CK(clk_i), .D(n_10120), .Q(u10_mem_b0_b_156), .SO(u10_mem_b0_b_156), .SE(scan_enable), .SI(u10_mem_b0_b_155));
SDFFNSRN u10_mem_reg_b0_b_b9_b (.CK(clk_i), .D(n_10118), .Q(u10_mem_b0_b_158), .SO(u10_mem_b0_b_158), .SE(scan_enable), .SI(u10_mem_b0_b_156));
SDFFN u10_wp_reg_b0_b (.CK(clk_i), .D(n_10333), .Q(n_9641), .SO(n_9641), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u10_mem_b0_b_158));
SDFFNSRN u11_din_tmp1_reg_b0_b (.CK(clk_i), .D(n_10115), .Q(u11_din_tmp1), .SO(u11_din_tmp1), .SE(scan_enable), .SI(n_9641));
SDFFNSRN u11_din_tmp1_reg_b10_b (.CK(clk_i), .D(n_10114), .Q(u11_din_tmp_51), .SO(u11_din_tmp_51), .SE(scan_enable), .SI(u11_din_tmp1));
SDFFNSRN u11_din_tmp1_reg_b11_b (.CK(clk_i), .D(n_10112), .Q(u11_din_tmp_52), .SO(u11_din_tmp_52), .SE(scan_enable), .SI(u11_din_tmp_51));
SDFFNSRN u11_din_tmp1_reg_b12_b (.CK(clk_i), .D(n_10111), .Q(u11_din_tmp_53), .SO(u11_din_tmp_53), .SE(scan_enable), .SI(u11_din_tmp_52));
SDFFNSRN u11_din_tmp1_reg_b13_b (.CK(clk_i), .D(n_10110), .Q(u11_din_tmp_54), .SO(u11_din_tmp_54), .SE(scan_enable), .SI(u11_din_tmp_53));
SDFFNSRN u11_din_tmp1_reg_b14_b (.CK(clk_i), .D(n_10108), .Q(u11_din_tmp_55), .SO(u11_din_tmp_55), .SE(scan_enable), .SI(u11_din_tmp_54));
SDFFNSRN u11_din_tmp1_reg_b15_b (.CK(clk_i), .D(n_10106), .Q(u11_din_tmp_56), .SO(u11_din_tmp_56), .SE(scan_enable), .SI(u11_din_tmp_55));
SDFFNSRN u11_din_tmp1_reg_b1_b (.CK(clk_i), .D(n_10105), .Q(u11_din_tmp_42), .SO(u11_din_tmp_42), .SE(scan_enable), .SI(u11_din_tmp_56));
SDFFNSRN u11_din_tmp1_reg_b2_b (.CK(clk_i), .D(n_10104), .Q(u11_din_tmp_43), .SO(u11_din_tmp_43), .SE(scan_enable), .SI(u11_din_tmp_42));
SDFFNSRN u11_din_tmp1_reg_b3_b (.CK(clk_i), .D(n_10102), .Q(u11_din_tmp_44), .SO(u11_din_tmp_44), .SE(scan_enable), .SI(u11_din_tmp_43));
SDFFNSRN u11_din_tmp1_reg_b5_b (.CK(clk_i), .D(n_10100), .Q(u11_din_tmp_46), .SO(u11_din_tmp_46), .SE(scan_enable), .SI(u11_din_tmp_44));
SDFFNSRN u11_din_tmp1_reg_b6_b (.CK(clk_i), .D(n_10099), .Q(u11_din_tmp_47), .SO(u11_din_tmp_47), .SE(scan_enable), .SI(u11_din_tmp_46));
SDFFNSRN u11_din_tmp1_reg_b7_b (.CK(clk_i), .D(n_10098), .Q(u11_din_tmp_48), .SO(u11_din_tmp_48), .SE(scan_enable), .SI(u11_din_tmp_47));
SDFFNSRN u11_din_tmp1_reg_b9_b (.CK(clk_i), .D(n_10096), .Q(u11_din_tmp_50), .SO(u11_din_tmp_50), .SE(scan_enable), .SI(u11_din_tmp_48));
SDFFNSRN u9_mem_reg_b2_b_b9_b (.CK(clk_i), .D(n_10264), .Q(u9_mem_b2_b_96), .SO(u9_mem_b2_b_96), .SE(scan_enable), .SI(u11_din_tmp_50));
SDFFN u18_int_set_reg_b1_b (.CK(clk_i), .D(n_10344), .Q(oc1_int_set_709), .SO(oc1_int_set_709), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u9_mem_b2_b_96));
SDFFN u19_int_set_reg_b1_b (.CK(clk_i), .D(n_10343), .Q(oc2_int_set_711), .SO(oc2_int_set_711), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc1_int_set_709));
SDFFN u24_int_set_reg_b2_b (.CK(clk_i), .D(n_10342), .Q(ic1_int_set_722), .SO(ic1_int_set_722), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc2_int_set_711));
SDFFN u15_crac_wr_reg (.CK(clk_i), .D(n_10339), .Q(crac_wr), .SO(crac_wr), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic1_int_set_722));
SDFFN u13_ints_r_reg_b1_b (.CK(clk_i), .D(n_10399), .Q(u13_ints_r_b1_b), .SO(u13_ints_r_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_wr));
SDFFNSRN u10_mem_reg_b0_b_b20_b (.CK(clk_i), .D(n_10130), .Q(u10_mem_b0_b_169), .SO(u10_mem_b0_b_169), .SE(scan_enable), .SI(u13_ints_r_b1_b));
SDFFNSRN u10_din_tmp1_reg_b13_b (.CK(clk_i), .D(n_9856), .Q(u10_din_tmp_54), .SO(u10_din_tmp_54), .SE(scan_enable), .SI(u10_mem_b0_b_169));
SDFFN u13_ints_r_reg_b26_b (.CK(clk_i), .D(n_10083), .Q(u13_ints_r_b26_b), .SO(u13_ints_r_b26_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u10_din_tmp_54));
SDFFNSRN u10_din_tmp1_reg_b11_b (.CK(clk_i), .D(n_9858), .Q(u10_din_tmp_52), .SO(u10_din_tmp_52), .SE(scan_enable), .SI(u13_ints_r_b26_b));
SDFFN u9_wp_reg_b0_b (.CK(clk_i), .D(n_9951), .Q(n_1203), .SO(n_1203), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u10_din_tmp_52));
SDFFNSRN u10_din_tmp1_reg_b5_b (.CK(clk_i), .D(n_9868), .Q(u10_din_tmp_46), .SO(u10_din_tmp_46), .SE(scan_enable), .SI(n_1203));
SDFFNSRN u10_din_tmp1_reg_b3_b (.CK(clk_i), .D(n_9871), .Q(u10_din_tmp_44), .SO(u10_din_tmp_44), .SE(scan_enable), .SI(u10_din_tmp_46));
SDFFNSRN u10_din_tmp1_reg_b1_b (.CK(clk_i), .D(n_9853), .Q(u10_din_tmp_42), .SO(u10_din_tmp_42), .SE(scan_enable), .SI(u10_din_tmp_44));
SDFFNSRN u10_din_tmp1_reg_b2_b (.CK(clk_i), .D(n_9872), .Q(u10_din_tmp_43), .SO(u10_din_tmp_43), .SE(scan_enable), .SI(u10_din_tmp_42));
SDFFNSRN u10_din_tmp1_reg_b4_b (.CK(clk_i), .D(n_9869), .Q(u10_din_tmp_45), .SO(u10_din_tmp_45), .SE(scan_enable), .SI(u10_din_tmp_43));
SDFFNSRN u10_din_tmp1_reg_b6_b (.CK(clk_i), .D(n_9867), .Q(u10_din_tmp_47), .SO(u10_din_tmp_47), .SE(scan_enable), .SI(u10_din_tmp_45));
SDFFNSRN u10_din_tmp1_reg_b8_b (.CK(clk_i), .D(n_9863), .Q(u10_din_tmp_49), .SO(u10_din_tmp_49), .SE(scan_enable), .SI(u10_din_tmp_47));
SDFFNSRN u10_din_tmp1_reg_b9_b (.CK(clk_i), .D(n_9862), .Q(u10_din_tmp_50), .SO(u10_din_tmp_50), .SE(scan_enable), .SI(u10_din_tmp_49));
SDFFNSRN u10_din_tmp1_reg_b7_b (.CK(clk_i), .D(n_9865), .Q(u10_din_tmp_48), .SO(u10_din_tmp_48), .SE(scan_enable), .SI(u10_din_tmp_50));
SDFFNSRN u10_din_tmp1_reg_b0_b (.CK(clk_i), .D(n_9861), .Q(u10_din_tmp1), .SO(u10_din_tmp1), .SE(scan_enable), .SI(u10_din_tmp_48));
SDFFNSRN u10_din_tmp1_reg_b10_b (.CK(clk_i), .D(n_9859), .Q(u10_din_tmp_51), .SO(u10_din_tmp_51), .SE(scan_enable), .SI(u10_din_tmp1));
SDFFNSRN u10_din_tmp1_reg_b15_b (.CK(clk_i), .D(n_9854), .Q(u10_din_tmp_56), .SO(u10_din_tmp_56), .SE(scan_enable), .SI(u10_din_tmp_51));
SDFFNSRN u10_din_tmp1_reg_b14_b (.CK(clk_i), .D(n_9855), .Q(u10_din_tmp_55), .SO(u10_din_tmp_55), .SE(scan_enable), .SI(u10_din_tmp_56));
SDFFNSRN u10_din_tmp1_reg_b12_b (.CK(clk_i), .D(n_9857), .Q(u10_din_tmp_53), .SO(u10_din_tmp_53), .SE(scan_enable), .SI(u10_din_tmp_55));
SDFFN u15_rdd1_reg (.CK(clk_i), .D(n_9884), .Q(u15_rdd1), .SO(u15_rdd1), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u10_din_tmp_53));
SDFFN u15_rdd2_reg (.CK(clk_i), .D(n_9883), .Q(u15_rdd2), .SO(u15_rdd2), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u15_rdd1));
SDFFN u20_int_set_reg_b0_b (.CK(clk_i), .D(n_10091), .Q(oc3_int_set), .SO(oc3_int_set), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u15_rdd2));
SDFFN u18_int_set_reg_b0_b (.CK(clk_i), .D(n_10092), .Q(oc1_int_set), .SO(oc1_int_set), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc3_int_set));
SDFFN u13_ints_r_reg_b23_b (.CK(clk_i), .D(n_9845), .Q(u13_ints_r_b23_b), .SO(u13_ints_r_b23_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc1_int_set));
SDFFN u13_ints_r_reg_b20_b (.CK(clk_i), .D(n_9846), .Q(u13_ints_r_b20_b), .SO(u13_ints_r_b20_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b23_b));
SDFFNSRN u9_wp_reg_b1_b (.CK(clk_i), .D(n_9836), .Q(u9_wp_b1_b), .SO(u9_wp_b1_b), .SE(scan_enable), .SI(u13_ints_r_b20_b));
SDFFNSRN u9_din_tmp1_reg_b9_b (.CK(clk_i), .D(n_9770), .Q(u9_din_tmp_50), .SO(u9_din_tmp_50), .SE(scan_enable), .SI(u9_wp_b1_b));
SDFFNSRN u9_din_tmp1_reg_b3_b (.CK(clk_i), .D(n_9776), .Q(u9_din_tmp_44), .SO(u9_din_tmp_44), .SE(scan_enable), .SI(u9_din_tmp_50));
SDFFNSRN u9_din_tmp1_reg_b10_b (.CK(clk_i), .D(n_9788), .Q(u9_din_tmp_51), .SO(u9_din_tmp_51), .SE(scan_enable), .SI(u9_din_tmp_44));
SDFFNSRN u9_din_tmp1_reg_b14_b (.CK(clk_i), .D(n_9782), .Q(u9_din_tmp_55), .SO(u9_din_tmp_55), .SE(scan_enable), .SI(u9_din_tmp_51));
SDFFNSRN u9_din_tmp1_reg_b0_b (.CK(clk_i), .D(n_9789), .Q(u9_din_tmp1), .SO(u9_din_tmp1), .SE(scan_enable), .SI(u9_din_tmp_55));
SDFFNSRN u9_din_tmp1_reg_b11_b (.CK(clk_i), .D(n_9786), .Q(u9_din_tmp_52), .SO(u9_din_tmp_52), .SE(scan_enable), .SI(u9_din_tmp1));
SDFFNSRN u9_din_tmp1_reg_b12_b (.CK(clk_i), .D(n_9785), .Q(u9_din_tmp_53), .SO(u9_din_tmp_53), .SE(scan_enable), .SI(u9_din_tmp_52));
SDFFNSRN u9_din_tmp1_reg_b13_b (.CK(clk_i), .D(n_9784), .Q(u9_din_tmp_54), .SO(u9_din_tmp_54), .SE(scan_enable), .SI(u9_din_tmp_53));
SDFFNSRN u9_din_tmp1_reg_b15_b (.CK(clk_i), .D(n_9780), .Q(u9_din_tmp_56), .SO(u9_din_tmp_56), .SE(scan_enable), .SI(u9_din_tmp_54));
SDFFNSRN u9_din_tmp1_reg_b1_b (.CK(clk_i), .D(n_9779), .Q(u9_din_tmp_42), .SO(u9_din_tmp_42), .SE(scan_enable), .SI(u9_din_tmp_56));
SDFFNSRN u9_din_tmp1_reg_b2_b (.CK(clk_i), .D(n_9778), .Q(u9_din_tmp_43), .SO(u9_din_tmp_43), .SE(scan_enable), .SI(u9_din_tmp_42));
SDFFNSRN u9_din_tmp1_reg_b5_b (.CK(clk_i), .D(n_9774), .Q(u9_din_tmp_46), .SO(u9_din_tmp_46), .SE(scan_enable), .SI(u9_din_tmp_43));
SDFFNSRN u9_din_tmp1_reg_b6_b (.CK(clk_i), .D(n_9773), .Q(u9_din_tmp_47), .SO(u9_din_tmp_47), .SE(scan_enable), .SI(u9_din_tmp_46));
SDFFNSRN u9_din_tmp1_reg_b4_b (.CK(clk_i), .D(n_9775), .Q(u9_din_tmp_45), .SO(u9_din_tmp_45), .SE(scan_enable), .SI(u9_din_tmp_47));
SDFFNSRN u9_din_tmp1_reg_b8_b (.CK(clk_i), .D(n_9771), .Q(u9_din_tmp_49), .SO(u9_din_tmp_49), .SE(scan_enable), .SI(u9_din_tmp_45));
SDFFNSRN u9_din_tmp1_reg_b7_b (.CK(clk_i), .D(n_9772), .Q(u9_din_tmp_48), .SO(u9_din_tmp_48), .SE(scan_enable), .SI(u9_din_tmp_49));
SDFFN u15_rdd3_reg (.CK(clk_i), .D(n_9796), .Q(u15_rdd3), .SO(u15_rdd3), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u9_din_tmp_48));
SDFFN u21_int_set_reg_b0_b (.CK(clk_i), .D(n_9848), .Q(oc4_int_set), .SO(oc4_int_set), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u15_rdd3));
SDFFN u22_int_set_reg_b0_b (.CK(clk_i), .D(n_9847), .Q(oc5_int_set), .SO(oc5_int_set), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc4_int_set));
SDFFN u17_int_set_reg_b0_b (.CK(clk_i), .D(n_9850), .Q(oc0_int_set), .SO(oc0_int_set), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc5_int_set));
SDFFN u19_int_set_reg_b0_b (.CK(clk_i), .D(n_9849), .Q(oc2_int_set), .SO(oc2_int_set), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc0_int_set));
SDFFNSRN u16_u8_dma_req_r1_reg (.CK(clk_i), .D(n_11907), .Q(u16_u8_dma_req_r1), .SO(u16_u8_dma_req_r1), .SE(scan_enable), .SI(oc2_int_set));
SDFFN u23_int_set_reg_b2_b (.CK(clk_i), .D(n_9758), .Q(ic0_int_set_720), .SO(ic0_int_set_720), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u16_u8_dma_req_r1));
SDFFNSRN u15_crac_rd_done_reg (.CK(clk_i), .D(n_9712), .Q(n_1036), .SO(n_1036), .SE(scan_enable), .SI(ic0_int_set_720));
SDFFNSRN u16_u6_dma_req_r1_reg (.CK(clk_i), .D(n_12374), .Q(n_12066), .SO(n_12066), .SE(scan_enable), .SI(n_1036));
SDFFNSRN u16_u7_dma_req_r1_reg (.CK(clk_i), .D(n_12379), .Q(n_12067), .SO(n_12067), .SE(scan_enable), .SI(n_12066));
SDFFN u14_u4_en_out_l_reg (.CK(clk_i), .D(n_9636), .Q(out_slt_18), .SO(out_slt_18), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(n_12067));
SDFFN u2_sync_resume_reg (.CK(clk_i), .D(n_9617), .Q(u2_sync_resume), .SO(u2_sync_resume), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(out_slt_18));
SDFFN u14_u0_en_out_l_reg (.CK(clk_i), .D(n_9640), .Q(out_slt_23), .SO(out_slt_23), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u2_sync_resume));
SDFFN u14_u1_en_out_l_reg (.CK(clk_i), .D(n_9639), .Q(out_slt_22), .SO(out_slt_22), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(out_slt_23));
SDFFN u14_u2_en_out_l_reg (.CK(clk_i), .D(n_9638), .Q(out_slt_20), .SO(out_slt_20), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(out_slt_22));
SDFFN u14_u3_en_out_l_reg (.CK(clk_i), .D(n_9637), .Q(out_slt_19), .SO(out_slt_19), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(out_slt_20));
SDFFN u14_u5_en_out_l_reg (.CK(clk_i), .D(n_9635), .Q(out_slt_17), .SO(out_slt_17), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(out_slt_19));
SDFFNSRN u14_crac_valid_r_reg (.CK(clk_i), .D(n_9629), .Q(out_slt_25), .SO(out_slt_25), .SE(scan_enable), .SI(out_slt_17));
SDFFN u26_ps_cnt_reg_b5_b (.CK(clk_i), .D(n_9593), .Q(u26_ps_cnt_b5_b), .SO(u26_ps_cnt_b5_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(out_slt_25));
SDFFN u26_ps_cnt_reg_b2_b (.CK(clk_i), .D(n_9596), .Q(n_760), .SO(n_760), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u26_ps_cnt_b5_b));
SDFFN u26_ps_cnt_reg_b0_b (.CK(clk_i), .D(n_9599), .Q(u26_ps_cnt_b0_b), .SO(u26_ps_cnt_b0_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(n_760));
SDFFN u26_ps_cnt_reg_b1_b (.CK(clk_i), .D(n_9598), .Q(u26_ps_cnt_b1_b), .SO(u26_ps_cnt_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u26_ps_cnt_b0_b));
SDFFN u26_ps_cnt_reg_b4_b (.CK(clk_i), .D(n_9594), .Q(u26_ps_cnt_b4_b), .SO(u26_ps_cnt_b4_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u26_ps_cnt_b1_b));
SDFFN u26_ps_cnt_reg_b3_b (.CK(clk_i), .D(n_9595), .Q(u26_ps_cnt_b3_b), .SO(u26_ps_cnt_b3_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u26_ps_cnt_b4_b));
SDFFNSRN u12_wb_data_o_reg_b1_b (.CK(clk_i), .D(n_9608), .Q(wb_data_o_b1_b), .SO(wb_data_o_b1_b), .SE(scan_enable), .SI(u26_ps_cnt_b3_b));
SDFFN u17_int_set_reg_b2_b (.CK(clk_i), .D(n_9578), .Q(oc0_int_set_708), .SO(oc0_int_set_708), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(wb_data_o_b1_b));
SDFFN u18_int_set_reg_b2_b (.CK(clk_i), .D(n_9577), .Q(oc1_int_set_710), .SO(oc1_int_set_710), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc0_int_set_708));
SDFFN u21_int_set_reg_b2_b (.CK(clk_i), .D(n_9574), .Q(oc4_int_set_716), .SO(oc4_int_set_716), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc1_int_set_710));
SDFFN u20_int_set_reg_b2_b (.CK(clk_i), .D(n_9575), .Q(oc3_int_set_714), .SO(oc3_int_set_714), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc4_int_set_716));
SDFFNSRN u14_crac_wr_r_reg (.CK(clk_i), .D(n_9580), .Q(out_slt_24), .SO(out_slt_24), .SE(scan_enable), .SI(oc3_int_set_714));
SDFFN u22_int_set_reg_b2_b (.CK(clk_i), .D(n_9573), .Q(oc5_int_set_718), .SO(oc5_int_set_718), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(out_slt_24));
SDFFN u19_int_set_reg_b2_b (.CK(clk_i), .D(n_9576), .Q(oc2_int_set_712), .SO(oc2_int_set_712), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc5_int_set_718));
SDFFNSRN u14_u3_full_empty_r_reg (.CK(clk_i), .D(n_9537), .Q(u14_u3_full_empty_r), .SO(u14_u3_full_empty_r), .SE(scan_enable), .SI(oc2_int_set_712));
SDFFN u25_int_set_reg_b0_b (.CK(clk_i), .D(n_9545), .Q(ic2_int_set), .SO(ic2_int_set), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u14_u3_full_empty_r));
SDFFNSRN u14_u0_full_empty_r_reg (.CK(clk_i), .D(n_9544), .Q(u14_u0_full_empty_r), .SO(u14_u0_full_empty_r), .SE(scan_enable), .SI(ic2_int_set));
SDFFNSRN u14_u1_full_empty_r_reg (.CK(clk_i), .D(n_9542), .Q(u14_u1_full_empty_r), .SO(u14_u1_full_empty_r), .SE(scan_enable), .SI(u14_u0_full_empty_r));
SDFFNSRN u14_u2_full_empty_r_reg (.CK(clk_i), .D(n_9539), .Q(u14_u2_full_empty_r), .SO(u14_u2_full_empty_r), .SE(scan_enable), .SI(u14_u1_full_empty_r));
SDFFNSRN u14_u5_full_empty_r_reg (.CK(clk_i), .D(n_9533), .Q(u14_u5_full_empty_r), .SO(u14_u5_full_empty_r), .SE(scan_enable), .SI(u14_u2_full_empty_r));
SDFFNSRN u14_u4_full_empty_r_reg (.CK(clk_i), .D(n_9535), .Q(u14_u4_full_empty_r), .SO(u14_u4_full_empty_r), .SE(scan_enable), .SI(u14_u5_full_empty_r));
SDFFNSRN u8_wp_reg_b0_b (.CK(clk_i), .D(n_9520), .Q(u8_wp_b0_b), .SO(u8_wp_b0_b), .SE(scan_enable), .SI(u14_u4_full_empty_r));
SDFFNSRN u3_wp_reg_b0_b (.CK(clk_i), .D(n_9519), .Q(u3_wp_b0_b), .SO(u3_wp_b0_b), .SE(scan_enable), .SI(u8_wp_b0_b));
SDFFNSRN u4_wp_reg_b0_b (.CK(clk_i), .D(n_9518), .Q(u4_wp_b0_b), .SO(u4_wp_b0_b), .SE(scan_enable), .SI(u3_wp_b0_b));
SDFFNSRN u5_wp_reg_b0_b (.CK(clk_i), .D(n_9517), .Q(u5_wp_b0_b), .SO(u5_wp_b0_b), .SE(scan_enable), .SI(u4_wp_b0_b));
SDFFNSRN u6_wp_reg_b0_b (.CK(clk_i), .D(n_9516), .Q(u6_wp_b0_b), .SO(u6_wp_b0_b), .SE(scan_enable), .SI(u5_wp_b0_b));
SDFFNSRN u7_wp_reg_b0_b (.CK(clk_i), .D(n_9515), .Q(u7_wp_b0_b), .SO(u7_wp_b0_b), .SE(scan_enable), .SI(u6_wp_b0_b));
SDFFN u26_ac97_rst__reg (.CK(clk_i), .D(n_9491), .Q(ac97_reset_pad_o_), .SO(ac97_reset_pad_o_), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_wp_b0_b));
SDFFN u26_cnt_reg_b2_b (.CK(clk_i), .D(n_9492), .Q(u26_cnt_b2_b), .SO(u26_cnt_b2_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ac97_reset_pad_o_));
SDFFN u23_int_set_reg_b0_b (.CK(clk_i), .D(n_9490), .Q(ic0_int_set), .SO(ic0_int_set), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u26_cnt_b2_b));
SDFFN u24_int_set_reg_b0_b (.CK(clk_i), .D(n_9485), .Q(ic1_int_set), .SO(ic1_int_set), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic0_int_set));
SDFFN u14_u8_en_out_l_reg (.CK(clk_i), .D(n_9461), .Q(u14_n_135), .SO(u14_n_135), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic1_int_set));
SDFFN u5_wp_reg_b1_b (.CK(clk_i), .D(n_9458), .Q(u5_wp_b1_b), .SO(u5_wp_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u14_n_135));
SDFFNSRN u6_wp_reg_b2_b (.CK(clk_i), .D(n_9465), .Q(u6_wp_b2_b), .SO(u6_wp_b2_b), .SE(scan_enable), .SI(u5_wp_b1_b));
SDFFN u26_cnt_reg_b0_b (.CK(clk_i), .D(n_9494), .Q(u26_cnt_b0_b), .SO(u26_cnt_b0_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_wp_b2_b));
SDFFN u26_cnt_reg_b1_b (.CK(clk_i), .D(n_9493), .Q(u26_cnt_b1_b), .SO(u26_cnt_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u26_cnt_b0_b));
SDFFNSRN u8_wp_reg_b2_b (.CK(clk_i), .D(n_9469), .Q(u8_wp_b2_b), .SO(u8_wp_b2_b), .SE(scan_enable), .SI(u26_cnt_b1_b));
SDFFNSRN u3_wp_reg_b2_b (.CK(clk_i), .D(n_9466), .Q(u3_wp_b2_b), .SO(u3_wp_b2_b), .SE(scan_enable), .SI(u8_wp_b2_b));
SDFFNSRN u5_wp_reg_b2_b (.CK(clk_i), .D(n_9467), .Q(u5_wp_b2_b), .SO(u5_wp_b2_b), .SE(scan_enable), .SI(u3_wp_b2_b));
SDFFNSRN u7_wp_reg_b2_b (.CK(clk_i), .D(n_9464), .Q(u7_wp_b2_b), .SO(u7_wp_b2_b), .SE(scan_enable), .SI(u5_wp_b2_b));
SDFFN u14_u6_en_out_l_reg (.CK(clk_i), .D(n_9463), .Q(u14_n_133), .SO(u14_n_133), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_wp_b2_b));
SDFFN u14_u7_en_out_l_reg (.CK(clk_i), .D(n_9462), .Q(u14_n_134), .SO(u14_n_134), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u14_n_133));
SDFFN u8_wp_reg_b1_b (.CK(clk_i), .D(n_9460), .Q(u8_wp_b1_b), .SO(u8_wp_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u14_n_134));
SDFFN u3_wp_reg_b1_b (.CK(clk_i), .D(n_9457), .Q(u3_wp_b1_b), .SO(u3_wp_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_wp_b1_b));
SDFFN u4_wp_reg_b1_b (.CK(clk_i), .D(n_9459), .Q(u4_wp_b1_b), .SO(u4_wp_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_wp_b1_b));
SDFFN u6_wp_reg_b1_b (.CK(clk_i), .D(n_9456), .Q(u6_wp_b1_b), .SO(u6_wp_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_wp_b1_b));
SDFFN u7_wp_reg_b1_b (.CK(clk_i), .D(n_9455), .Q(u7_wp_b1_b), .SO(u7_wp_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_wp_b1_b));
SDFFNSRN u4_wp_reg_b2_b (.CK(clk_i), .D(n_9468), .Q(u4_wp_b2_b), .SO(u4_wp_b2_b), .SE(scan_enable), .SI(u7_wp_b1_b));
SDFFNSRN u15_valid_r_reg (.CK(clk_i), .D(n_11823), .Q(u15_valid_r), .SO(u15_valid_r), .SE(scan_enable), .SI(u4_wp_b2_b));
SDFFN u4_mem_reg_b0_b_b13_b (.CK(clk_i), .D(n_9442), .Q(u4_mem_b0_b_103), .SO(u4_mem_b0_b_103), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u15_valid_r));
SDFFN u4_mem_reg_b0_b_b14_b (.CK(clk_i), .D(n_9441), .Q(u4_mem_b0_b_104), .SO(u4_mem_b0_b_104), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_103));
SDFFN u4_mem_reg_b0_b_b16_b (.CK(clk_i), .D(n_9440), .Q(u4_mem_b0_b_106), .SO(u4_mem_b0_b_106), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_104));
SDFFN u4_mem_reg_b0_b_b19_b (.CK(clk_i), .D(n_9439), .Q(u4_mem_b0_b_109), .SO(u4_mem_b0_b_109), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_106));
SDFFN u4_mem_reg_b0_b_b22_b (.CK(clk_i), .D(n_9437), .Q(u4_mem_b0_b_112), .SO(u4_mem_b0_b_112), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_109));
SDFFN u4_mem_reg_b0_b_b24_b (.CK(clk_i), .D(n_9435), .Q(u4_mem_b0_b_114), .SO(u4_mem_b0_b_114), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_112));
SDFFN u4_mem_reg_b0_b_b31_b (.CK(clk_i), .D(n_9434), .Q(u4_mem_b0_b_121), .SO(u4_mem_b0_b_121), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_114));
SDFFN u4_mem_reg_b0_b_b4_b (.CK(clk_i), .D(n_9433), .Q(u4_mem_b0_b_94), .SO(u4_mem_b0_b_94), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_121));
SDFFN u4_mem_reg_b0_b_b7_b (.CK(clk_i), .D(n_9432), .Q(u4_mem_b0_b_97), .SO(u4_mem_b0_b_97), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_94));
SDFFN u4_mem_reg_b0_b_b9_b (.CK(clk_i), .D(n_9430), .Q(u4_mem_b0_b_99), .SO(u4_mem_b0_b_99), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_97));
SDFFN u5_mem_reg_b0_b_b13_b (.CK(clk_i), .D(n_9429), .Q(u5_mem_b0_b_103), .SO(u5_mem_b0_b_103), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_99));
SDFFN u5_mem_reg_b0_b_b14_b (.CK(clk_i), .D(n_9428), .Q(u5_mem_b0_b_104), .SO(u5_mem_b0_b_104), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_103));
SDFFN u5_mem_reg_b0_b_b16_b (.CK(clk_i), .D(n_9427), .Q(u5_mem_b0_b_106), .SO(u5_mem_b0_b_106), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_104));
SDFFN u5_mem_reg_b0_b_b19_b (.CK(clk_i), .D(n_9426), .Q(u5_mem_b0_b_109), .SO(u5_mem_b0_b_109), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_106));
SDFFN u5_mem_reg_b0_b_b22_b (.CK(clk_i), .D(n_9424), .Q(u5_mem_b0_b_112), .SO(u5_mem_b0_b_112), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_109));
SDFFN u5_mem_reg_b0_b_b24_b (.CK(clk_i), .D(n_9422), .Q(u5_mem_b0_b_114), .SO(u5_mem_b0_b_114), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_112));
SDFFN u5_mem_reg_b0_b_b31_b (.CK(clk_i), .D(n_9421), .Q(u5_mem_b0_b_121), .SO(u5_mem_b0_b_121), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_114));
SDFFN u5_mem_reg_b0_b_b4_b (.CK(clk_i), .D(n_9420), .Q(u5_mem_b0_b_94), .SO(u5_mem_b0_b_94), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_121));
SDFFN u5_mem_reg_b0_b_b7_b (.CK(clk_i), .D(n_9419), .Q(u5_mem_b0_b_97), .SO(u5_mem_b0_b_97), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_94));
SDFFN u5_mem_reg_b0_b_b9_b (.CK(clk_i), .D(n_9417), .Q(u5_mem_b0_b_99), .SO(u5_mem_b0_b_99), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_97));
SDFFN u6_mem_reg_b0_b_b13_b (.CK(clk_i), .D(n_9414), .Q(u6_mem_b0_b_103), .SO(u6_mem_b0_b_103), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_99));
SDFFN u6_mem_reg_b0_b_b14_b (.CK(clk_i), .D(n_9413), .Q(u6_mem_b0_b_104), .SO(u6_mem_b0_b_104), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_103));
SDFFN u6_mem_reg_b0_b_b16_b (.CK(clk_i), .D(n_9412), .Q(u6_mem_b0_b_106), .SO(u6_mem_b0_b_106), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_104));
SDFFN u6_mem_reg_b0_b_b19_b (.CK(clk_i), .D(n_9411), .Q(u6_mem_b0_b_109), .SO(u6_mem_b0_b_109), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_106));
SDFFN u6_mem_reg_b0_b_b22_b (.CK(clk_i), .D(n_9409), .Q(u6_mem_b0_b_112), .SO(u6_mem_b0_b_112), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_109));
SDFFN u6_mem_reg_b0_b_b24_b (.CK(clk_i), .D(n_9407), .Q(u6_mem_b0_b_114), .SO(u6_mem_b0_b_114), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_112));
SDFFN u6_mem_reg_b0_b_b31_b (.CK(clk_i), .D(n_9406), .Q(u6_mem_b0_b_121), .SO(u6_mem_b0_b_121), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_114));
SDFFN u6_mem_reg_b0_b_b4_b (.CK(clk_i), .D(n_9405), .Q(u6_mem_b0_b_94), .SO(u6_mem_b0_b_94), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_121));
SDFFN u6_mem_reg_b0_b_b7_b (.CK(clk_i), .D(n_9404), .Q(u6_mem_b0_b_97), .SO(u6_mem_b0_b_97), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_94));
SDFFN u6_mem_reg_b0_b_b9_b (.CK(clk_i), .D(n_9402), .Q(u6_mem_b0_b_99), .SO(u6_mem_b0_b_99), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_97));
SDFFN u7_mem_reg_b0_b_b13_b (.CK(clk_i), .D(n_9401), .Q(u7_mem_b0_b_103), .SO(u7_mem_b0_b_103), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_99));
SDFFN u7_mem_reg_b0_b_b14_b (.CK(clk_i), .D(n_9400), .Q(u7_mem_b0_b_104), .SO(u7_mem_b0_b_104), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_103));
SDFFN u7_mem_reg_b0_b_b16_b (.CK(clk_i), .D(n_9399), .Q(u7_mem_b0_b_106), .SO(u7_mem_b0_b_106), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_104));
SDFFN u7_mem_reg_b0_b_b19_b (.CK(clk_i), .D(n_9398), .Q(u7_mem_b0_b_109), .SO(u7_mem_b0_b_109), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_106));
SDFFN u7_mem_reg_b0_b_b22_b (.CK(clk_i), .D(n_9396), .Q(u7_mem_b0_b_112), .SO(u7_mem_b0_b_112), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_109));
SDFFN u7_mem_reg_b0_b_b24_b (.CK(clk_i), .D(n_9394), .Q(u7_mem_b0_b_114), .SO(u7_mem_b0_b_114), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_112));
SDFFN u7_mem_reg_b0_b_b31_b (.CK(clk_i), .D(n_9393), .Q(u7_mem_b0_b_121), .SO(u7_mem_b0_b_121), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_114));
SDFFN u7_mem_reg_b0_b_b4_b (.CK(clk_i), .D(n_9392), .Q(u7_mem_b0_b_94), .SO(u7_mem_b0_b_94), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_121));
SDFFN u7_mem_reg_b0_b_b7_b (.CK(clk_i), .D(n_9391), .Q(u7_mem_b0_b_97), .SO(u7_mem_b0_b_97), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_94));
SDFFN u7_mem_reg_b0_b_b9_b (.CK(clk_i), .D(n_9389), .Q(u7_mem_b0_b_99), .SO(u7_mem_b0_b_99), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_97));
SDFFN u3_mem_reg_b0_b_b11_b (.CK(clk_i), .D(n_9443), .Q(u3_mem_b0_b_101), .SO(u3_mem_b0_b_101), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_99));
SDFFN u3_mem_reg_b0_b_b12_b (.CK(clk_i), .D(n_9388), .Q(u3_mem_b0_b_102), .SO(u3_mem_b0_b_102), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_101));
SDFFN u3_mem_reg_b0_b_b15_b (.CK(clk_i), .D(n_9387), .Q(u3_mem_b0_b_105), .SO(u3_mem_b0_b_105), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_102));
SDFFN u8_mem_reg_b0_b_b0_b (.CK(clk_i), .D(n_9386), .Q(u8_mem_b0_b), .SO(u8_mem_b0_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_105));
SDFFN u8_mem_reg_b0_b_b11_b (.CK(clk_i), .D(n_9385), .Q(u8_mem_b0_b_101), .SO(u8_mem_b0_b_101), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b));
SDFFN u8_mem_reg_b0_b_b12_b (.CK(clk_i), .D(n_9383), .Q(u8_mem_b0_b_102), .SO(u8_mem_b0_b_102), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_101));
SDFFN u8_mem_reg_b0_b_b17_b (.CK(clk_i), .D(n_9381), .Q(u8_mem_b0_b_107), .SO(u8_mem_b0_b_107), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_102));
SDFFN u3_mem_reg_b0_b_b1_b (.CK(clk_i), .D(n_9382), .Q(u3_mem_b0_b_91), .SO(u3_mem_b0_b_91), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_107));
SDFFN u3_mem_reg_b0_b_b21_b (.CK(clk_i), .D(n_9380), .Q(u3_mem_b0_b_111), .SO(u3_mem_b0_b_111), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_91));
SDFFN u8_mem_reg_b0_b_b26_b (.CK(clk_i), .D(n_9379), .Q(u8_mem_b0_b_116), .SO(u8_mem_b0_b_116), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_111));
SDFFN u8_mem_reg_b0_b_b28_b (.CK(clk_i), .D(n_9378), .Q(u8_mem_b0_b_118), .SO(u8_mem_b0_b_118), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_116));
SDFFN u8_mem_reg_b0_b_b29_b (.CK(clk_i), .D(n_9376), .Q(u8_mem_b0_b_119), .SO(u8_mem_b0_b_119), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_118));
SDFFN u8_mem_reg_b0_b_b30_b (.CK(clk_i), .D(n_9375), .Q(u8_mem_b0_b_120), .SO(u8_mem_b0_b_120), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_119));
SDFFN u3_mem_reg_b0_b_b27_b (.CK(clk_i), .D(n_9373), .Q(u3_mem_b0_b_117), .SO(u3_mem_b0_b_117), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_120));
SDFFN u8_mem_reg_b0_b_b4_b (.CK(clk_i), .D(n_9371), .Q(u8_mem_b0_b_94), .SO(u8_mem_b0_b_94), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_117));
SDFFN u8_mem_reg_b0_b_b5_b (.CK(clk_i), .D(n_9370), .Q(u8_mem_b0_b_95), .SO(u8_mem_b0_b_95), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_94));
SDFFN u3_mem_reg_b0_b_b2_b (.CK(clk_i), .D(n_9416), .Q(u3_mem_b0_b_92), .SO(u3_mem_b0_b_92), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_95));
SDFFN u3_mem_reg_b0_b_b29_b (.CK(clk_i), .D(n_9369), .Q(u3_mem_b0_b_119), .SO(u3_mem_b0_b_119), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_92));
SDFFN u3_mem_reg_b0_b_b6_b (.CK(clk_i), .D(n_9366), .Q(u3_mem_b0_b_96), .SO(u3_mem_b0_b_96), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_119));
SDFFN u3_mem_reg_b0_b_b5_b (.CK(clk_i), .D(n_9368), .Q(u3_mem_b0_b_95), .SO(u3_mem_b0_b_95), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_96));
SDFFN u13_crac_r_reg_b6_b (.CK(clk_i), .D(n_8627), .Q(crac_out_867), .SO(crac_out_867), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_95));
SDFFN u3_mem_reg_b0_b_b17_b (.CK(clk_i), .D(n_8720), .Q(u3_mem_b0_b_107), .SO(u3_mem_b0_b_107), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_out_867));
SDFFN u8_mem_reg_b2_b_b18_b (.CK(clk_i), .D(n_8875), .Q(u8_mem_b2_b_46), .SO(u8_mem_b2_b_46), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_107));
SDFFN u7_mem_reg_b0_b_b20_b (.CK(clk_i), .D(n_8742), .Q(u7_mem_b0_b_110), .SO(u7_mem_b0_b_110), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_46));
SDFFN u8_mem_reg_b2_b_b25_b (.CK(clk_i), .D(n_8861), .Q(u8_mem_b2_b_53), .SO(u8_mem_b2_b_53), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_110));
SDFFN u8_mem_reg_b2_b_b28_b (.CK(clk_i), .D(n_8855), .Q(u8_mem_b2_b_56), .SO(u8_mem_b2_b_56), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_53));
SDFFN u4_mem_reg_b2_b_b16_b (.CK(clk_i), .D(n_8294), .Q(u4_mem_b2_b_44), .SO(u4_mem_b2_b_44), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_56));
SDFFN u5_mem_reg_b1_b_b26_b (.CK(clk_i), .D(n_9293), .Q(u5_mem_b1_b_85), .SO(u5_mem_b1_b_85), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_44));
SDFFN u13_occ0_r_reg_b11_b (.CK(clk_i), .D(n_8569), .Q(oc1_cfg_976), .SO(oc1_cfg_976), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_85));
SDFFN u5_mem_reg_b1_b_b22_b (.CK(clk_i), .D(n_9298), .Q(u5_mem_b1_b_81), .SO(u5_mem_b1_b_81), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc1_cfg_976));
SDFFN u5_mem_reg_b1_b_b15_b (.CK(clk_i), .D(n_9310), .Q(u5_mem_b1_b_74), .SO(u5_mem_b1_b_74), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_81));
SDFFN u5_mem_reg_b1_b_b19_b (.CK(clk_i), .D(n_9302), .Q(u5_mem_b1_b_78), .SO(u5_mem_b1_b_78), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_74));
SDFFN u5_mem_reg_b1_b_b11_b (.CK(clk_i), .D(n_9315), .Q(u5_mem_b1_b_70), .SO(u5_mem_b1_b_70), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_78));
SDFFN u3_mem_reg_b1_b_b22_b (.CK(clk_i), .D(n_8866), .Q(u3_mem_b1_b_81), .SO(u3_mem_b1_b_81), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_70));
SDFFN u8_mem_reg_b2_b_b20_b (.CK(clk_i), .D(n_8869), .Q(u8_mem_b2_b_48), .SO(u8_mem_b2_b_48), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_81));
SDFFN u4_mem_reg_b3_b_b9_b (.CK(clk_i), .D(n_9319), .Q(u4_mem_b3_b_130), .SO(u4_mem_b3_b_130), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_48));
SDFFN u4_mem_reg_b3_b_b5_b (.CK(clk_i), .D(n_9324), .Q(u4_mem_b3_b_126), .SO(u4_mem_b3_b_126), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_130));
SDFFN u4_mem_reg_b3_b_b30_b (.CK(clk_i), .D(n_9329), .Q(u4_mem_b3_b_151), .SO(u4_mem_b3_b_151), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_126));
SDFFN u8_mem_reg_b0_b_b15_b (.CK(clk_i), .D(n_8715), .Q(u8_mem_b0_b_105), .SO(u8_mem_b0_b_105), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_151));
SDFFN u3_mem_reg_b0_b_b16_b (.CK(clk_i), .D(n_8722), .Q(u3_mem_b0_b_106), .SO(u3_mem_b0_b_106), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_105));
SDFFN u4_mem_reg_b3_b_b23_b (.CK(clk_i), .D(n_9339), .Q(u4_mem_b3_b_144), .SO(u4_mem_b3_b_144), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_106));
SDFFN u4_mem_reg_b3_b_b27_b (.CK(clk_i), .D(n_9334), .Q(u4_mem_b3_b_148), .SO(u4_mem_b3_b_148), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_144));
SDFFN u8_mem_reg_b1_b_b6_b (.CK(clk_i), .D(n_9072), .Q(u8_mem_b1_b_65), .SO(u8_mem_b1_b_65), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_148));
SDFFN u13_occ0_r_reg_b8_b (.CK(clk_i), .D(n_8523), .Q(oc1_cfg), .SO(oc1_cfg), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_65));
SDFFN u13_icc_r_reg_b8_b (.CK(clk_i), .D(n_8575), .Q(ic1_cfg), .SO(ic1_cfg), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc1_cfg));
SDFFN u8_mem_reg_b2_b_b13_b (.CK(clk_i), .D(n_8882), .Q(u8_mem_b2_b_41), .SO(u8_mem_b2_b_41), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic1_cfg));
SDFFN u3_mem_reg_b1_b_b19_b (.CK(clk_i), .D(n_8880), .Q(u3_mem_b1_b_78), .SO(u3_mem_b1_b_78), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_41));
SDFFN u4_mem_reg_b2_b_b9_b (.CK(clk_i), .D(n_8266), .Q(u4_mem_b2_b_37), .SO(u4_mem_b2_b_37), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_78));
SDFFN u4_mem_reg_b3_b_b16_b (.CK(clk_i), .D(n_9350), .Q(u4_mem_b3_b_137), .SO(u4_mem_b3_b_137), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_37));
SDFFN u4_mem_reg_b3_b_b12_b (.CK(clk_i), .D(n_8261), .Q(u4_mem_b3_b_133), .SO(u4_mem_b3_b_133), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_137));
SDFFN u4_mem_reg_b2_b_b5_b (.CK(clk_i), .D(n_8270), .Q(u4_mem_b2_b_33), .SO(u4_mem_b2_b_33), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_133));
SDFFN u3_mem_reg_b1_b_b15_b (.CK(clk_i), .D(n_8897), .Q(u3_mem_b1_b_74), .SO(u3_mem_b1_b_74), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_33));
SDFFN u4_mem_reg_b2_b_b30_b (.CK(clk_i), .D(n_8274), .Q(u4_mem_b2_b_58), .SO(u4_mem_b2_b_58), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_74));
SDFFN u4_mem_reg_b2_b_b27_b (.CK(clk_i), .D(n_8280), .Q(u4_mem_b2_b_55), .SO(u4_mem_b2_b_55), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_58));
SDFFN u4_mem_reg_b2_b_b23_b (.CK(clk_i), .D(n_8284), .Q(u4_mem_b2_b_51), .SO(u4_mem_b2_b_51), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_55));
SDFFN u7_mem_reg_b0_b_b30_b (.CK(clk_i), .D(n_8731), .Q(u7_mem_b0_b_120), .SO(u7_mem_b0_b_120), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_51));
SDFFN u3_mem_reg_b2_b_b2_b (.CK(clk_i), .D(n_8400), .Q(u3_mem_b2_b_30), .SO(u3_mem_b2_b_30), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_120));
SDFFN u8_mem_reg_b1_b_b21_b (.CK(clk_i), .D(n_8924), .Q(u8_mem_b1_b_80), .SO(u8_mem_b1_b_80), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_30));
SDFFN u3_mem_reg_b1_b_b11_b (.CK(clk_i), .D(n_8908), .Q(u3_mem_b1_b_70), .SO(u3_mem_b1_b_70), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_80));
SDFFN u8_mem_reg_b1_b_b3_b (.CK(clk_i), .D(n_8902), .Q(u8_mem_b1_b_62), .SO(u8_mem_b1_b_62), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_70));
SDFFN u4_mem_reg_b2_b_b12_b (.CK(clk_i), .D(n_8298), .Q(u4_mem_b2_b_40), .SO(u4_mem_b2_b_40), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_62));
SDFFN u4_mem_reg_b1_b_b30_b (.CK(clk_i), .D(n_8313), .Q(u4_mem_b1_b_89), .SO(u4_mem_b1_b_89), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_40));
SDFFN u4_mem_reg_b1_b_b9_b (.CK(clk_i), .D(n_8303), .Q(u4_mem_b1_b_68), .SO(u4_mem_b1_b_68), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_89));
SDFFN u4_mem_reg_b1_b_b5_b (.CK(clk_i), .D(n_8308), .Q(u4_mem_b1_b_64), .SO(u4_mem_b1_b_64), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_68));
SDFFN u4_mem_reg_b1_b_b27_b (.CK(clk_i), .D(n_8320), .Q(u4_mem_b1_b_86), .SO(u4_mem_b1_b_86), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_64));
SDFFN u8_mem_reg_b1_b_b28_b (.CK(clk_i), .D(n_9196), .Q(u8_mem_b1_b_87), .SO(u8_mem_b1_b_87), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_86));
SDFFN u3_mem_reg_b0_b_b13_b (.CK(clk_i), .D(n_8724), .Q(u3_mem_b0_b_103), .SO(u3_mem_b0_b_103), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_87));
SDFFN u8_mem_reg_b1_b_b25_b (.CK(clk_i), .D(n_8918), .Q(u8_mem_b1_b_84), .SO(u8_mem_b1_b_84), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_103));
SDFFN u4_mem_reg_b1_b_b23_b (.CK(clk_i), .D(n_8325), .Q(u4_mem_b1_b_82), .SO(u4_mem_b1_b_82), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_84));
SDFFN u4_mem_reg_b1_b_b16_b (.CK(clk_i), .D(n_8336), .Q(u4_mem_b1_b_75), .SO(u4_mem_b1_b_75), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_82));
SDFFN u7_mem_reg_b0_b_b6_b (.CK(clk_i), .D(n_8727), .Q(u7_mem_b0_b_96), .SO(u7_mem_b0_b_96), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_75));
SDFFN u7_mem_reg_b1_b_b25_b (.CK(clk_i), .D(n_9042), .Q(u7_mem_b1_b_84), .SO(u7_mem_b1_b_84), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_96));
SDFFN u3_mem_reg_b3_b_b3_b (.CK(clk_i), .D(n_9069), .Q(u3_mem_b3_b_124), .SO(u3_mem_b3_b_124), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_84));
SDFFN u4_mem_reg_b1_b_b12_b (.CK(clk_i), .D(n_8342), .Q(u4_mem_b1_b_71), .SO(u4_mem_b1_b_71), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_124));
SDFFN u7_mem_reg_b3_b_b3_b (.CK(clk_i), .D(n_8952), .Q(u7_mem_b3_b_124), .SO(u7_mem_b3_b_124), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_71));
SDFFN u8_mem_reg_b1_b_b14_b (.CK(clk_i), .D(n_8935), .Q(u8_mem_b1_b_73), .SO(u8_mem_b1_b_73), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_124));
SDFFN u8_mem_reg_b1_b_b18_b (.CK(clk_i), .D(n_8929), .Q(u8_mem_b1_b_77), .SO(u8_mem_b1_b_77), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_73));
SDFFN u3_mem_reg_b3_b_b6_b (.CK(clk_i), .D(n_8355), .Q(u3_mem_b3_b_127), .SO(u3_mem_b3_b_127), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_77));
SDFFN u3_mem_reg_b3_b_b22_b (.CK(clk_i), .D(n_8371), .Q(u3_mem_b3_b_143), .SO(u3_mem_b3_b_143), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_127));
SDFFN u3_mem_reg_b3_b_b30_b (.CK(clk_i), .D(n_8361), .Q(u3_mem_b3_b_151), .SO(u3_mem_b3_b_151), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_143));
SDFFN u3_mem_reg_b3_b_b27_b (.CK(clk_i), .D(n_8366), .Q(u3_mem_b3_b_148), .SO(u3_mem_b3_b_148), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_151));
SDFFN u7_mem_reg_b0_b_b23_b (.CK(clk_i), .D(n_8739), .Q(u7_mem_b0_b_113), .SO(u7_mem_b0_b_113), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_148));
SDFFN u3_mem_reg_b3_b_b19_b (.CK(clk_i), .D(n_8376), .Q(u3_mem_b3_b_140), .SO(u3_mem_b3_b_140), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_113));
SDFFNSRN u14_u0_en_out_l2_reg (.CK(clk_i), .D(n_9480), .Q(n_11507), .SO(n_11507), .SE(scan_enable), .SI(u3_mem_b3_b_140));
SDFFNSRN u14_u1_en_out_l2_reg (.CK(clk_i), .D(n_9479), .Q(u14_u1_en_out_l2), .SO(u14_u1_en_out_l2), .SE(scan_enable), .SI(n_11507));
SDFFNSRN u14_u2_en_out_l2_reg (.CK(clk_i), .D(n_9478), .Q(n_11533), .SO(n_11533), .SE(scan_enable), .SI(u14_u1_en_out_l2));
SDFFNSRN u14_u3_en_out_l2_reg (.CK(clk_i), .D(n_9477), .Q(n_11529), .SO(n_11529), .SE(scan_enable), .SI(n_11533));
SDFFNSRN u14_u4_en_out_l2_reg (.CK(clk_i), .D(n_9476), .Q(n_11528), .SO(n_11528), .SE(scan_enable), .SI(n_11529));
SDFFNSRN u14_u5_en_out_l2_reg (.CK(clk_i), .D(n_9475), .Q(n_11530), .SO(n_11530), .SE(scan_enable), .SI(n_11528));
SDFFN u6_mem_reg_b0_b_b12_b (.CK(clk_i), .D(n_8778), .Q(u6_mem_b0_b_102), .SO(u6_mem_b0_b_102), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(n_11530));
SDFFN u8_mem_reg_b1_b_b10_b (.CK(clk_i), .D(n_8940), .Q(u8_mem_b1_b_69), .SO(u8_mem_b1_b_69), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_102));
SDFFN u7_mem_reg_b3_b_b7_b (.CK(clk_i), .D(n_8946), .Q(u7_mem_b3_b_128), .SO(u7_mem_b3_b_128), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_69));
SDFFN u3_mem_reg_b3_b_b15_b (.CK(clk_i), .D(n_8381), .Q(u3_mem_b3_b_136), .SO(u3_mem_b3_b_136), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_128));
SDFFN u3_mem_reg_b3_b_b11_b (.CK(clk_i), .D(n_8386), .Q(u3_mem_b3_b_132), .SO(u3_mem_b3_b_132), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_136));
SDFFN u3_mem_reg_b2_b_b8_b (.CK(clk_i), .D(n_8391), .Q(u3_mem_b2_b_36), .SO(u3_mem_b2_b_36), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_132));
SDFFN u7_mem_reg_b0_b_b12_b (.CK(clk_i), .D(n_8750), .Q(u7_mem_b0_b_102), .SO(u7_mem_b0_b_102), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_36));
SDFFN u7_mem_reg_b3_b_b14_b (.CK(clk_i), .D(n_8977), .Q(u7_mem_b3_b_135), .SO(u7_mem_b3_b_135), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_102));
SDFFN u7_mem_reg_b3_b_b25_b (.CK(clk_i), .D(n_8962), .Q(u7_mem_b3_b_146), .SO(u7_mem_b3_b_146), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_135));
SDFFN u7_mem_reg_b3_b_b29_b (.CK(clk_i), .D(n_8956), .Q(u7_mem_b3_b_150), .SO(u7_mem_b3_b_150), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_146));
SDFFN u3_mem_reg_b2_b_b26_b (.CK(clk_i), .D(n_8404), .Q(u3_mem_b2_b_54), .SO(u3_mem_b2_b_54), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_150));
SDFFN u3_mem_reg_b2_b_b22_b (.CK(clk_i), .D(n_8406), .Q(u3_mem_b2_b_50), .SO(u3_mem_b2_b_50), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_54));
SDFFN u3_mem_reg_b2_b_b18_b (.CK(clk_i), .D(n_8412), .Q(u3_mem_b2_b_46), .SO(u3_mem_b2_b_46), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_50));
SDFFN u8_mem_reg_b3_b_b8_b (.CK(clk_i), .D(n_9068), .Q(u8_mem_b3_b_129), .SO(u8_mem_b3_b_129), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_46));
SDFFN u8_mem_reg_b3_b_b6_b (.CK(clk_i), .D(n_9197), .Q(u8_mem_b3_b_127), .SO(u8_mem_b3_b_127), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_129));
SDFFN u7_mem_reg_b3_b_b21_b (.CK(clk_i), .D(n_8967), .Q(u7_mem_b3_b_142), .SO(u7_mem_b3_b_142), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_127));
SDFFN u7_mem_reg_b3_b_b18_b (.CK(clk_i), .D(n_8972), .Q(u7_mem_b3_b_139), .SO(u7_mem_b3_b_139), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_142));
SDFFN u8_mem_reg_b3_b_b3_b (.CK(clk_i), .D(n_8422), .Q(u8_mem_b3_b_124), .SO(u8_mem_b3_b_124), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_139));
SDFFN u3_mem_reg_b2_b_b11_b (.CK(clk_i), .D(n_8427), .Q(u3_mem_b2_b_39), .SO(u3_mem_b2_b_39), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_124));
SDFFN u8_mem_reg_b3_b_b28_b (.CK(clk_i), .D(n_8365), .Q(u8_mem_b3_b_149), .SO(u8_mem_b3_b_149), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_39));
SDFFN u7_mem_reg_b0_b_b17_b (.CK(clk_i), .D(n_8747), .Q(u7_mem_b0_b_107), .SO(u7_mem_b0_b_107), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_149));
SDFFN u7_mem_reg_b0_b_b0_b (.CK(clk_i), .D(n_8753), .Q(u7_mem_b0_b), .SO(u7_mem_b0_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_107));
SDFFN u8_mem_reg_b3_b_b22_b (.CK(clk_i), .D(n_8439), .Q(u8_mem_b3_b_143), .SO(u8_mem_b3_b_143), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b));
SDFFN u8_mem_reg_b3_b_b25_b (.CK(clk_i), .D(n_8434), .Q(u8_mem_b3_b_146), .SO(u8_mem_b3_b_146), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_143));
SDFFN u7_mem_reg_b2_b_b25_b (.CK(clk_i), .D(n_9000), .Q(u7_mem_b2_b_53), .SO(u7_mem_b2_b_53), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_146));
SDFFN u7_mem_reg_b2_b_b7_b (.CK(clk_i), .D(n_8986), .Q(u7_mem_b2_b_35), .SO(u7_mem_b2_b_35), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_53));
SDFFN u7_mem_reg_b3_b_b10_b (.CK(clk_i), .D(n_8982), .Q(u7_mem_b3_b_131), .SO(u7_mem_b3_b_131), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_35));
SDFFN u8_mem_reg_b3_b_b18_b (.CK(clk_i), .D(n_8448), .Q(u8_mem_b3_b_139), .SO(u8_mem_b3_b_139), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_131));
SDFFN u3_mem_reg_b1_b_b3_b (.CK(clk_i), .D(n_8460), .Q(u3_mem_b1_b_62), .SO(u3_mem_b1_b_62), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_139));
SDFFN u8_mem_reg_b3_b_b15_b (.CK(clk_i), .D(n_8456), .Q(u8_mem_b3_b_136), .SO(u8_mem_b3_b_136), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_62));
SDFFN u8_mem_reg_b3_b_b10_b (.CK(clk_i), .D(n_8465), .Q(u8_mem_b3_b_131), .SO(u8_mem_b3_b_131), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_136));
SDFFN u7_mem_reg_b2_b_b3_b (.CK(clk_i), .D(n_8990), .Q(u7_mem_b2_b_31), .SO(u7_mem_b2_b_31), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_131));
SDFFN u7_mem_reg_b2_b_b29_b (.CK(clk_i), .D(n_8995), .Q(u7_mem_b2_b_57), .SO(u7_mem_b2_b_57), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_31));
SDFFN u3_mem_reg_b1_b_b2_b (.CK(clk_i), .D(n_8471), .Q(u3_mem_b1_b_61), .SO(u3_mem_b1_b_61), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_57));
SDFFN u7_mem_reg_b2_b_b21_b (.CK(clk_i), .D(n_9004), .Q(u7_mem_b2_b_49), .SO(u7_mem_b2_b_49), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_61));
SDFFN u7_mem_reg_b2_b_b18_b (.CK(clk_i), .D(n_9009), .Q(u7_mem_b2_b_46), .SO(u7_mem_b2_b_46), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_49));
SDFFN u6_mem_reg_b0_b_b30_b (.CK(clk_i), .D(n_8759), .Q(u6_mem_b0_b_120), .SO(u6_mem_b0_b_120), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_46));
SDFFN u6_mem_reg_b0_b_b6_b (.CK(clk_i), .D(n_8755), .Q(u6_mem_b0_b_96), .SO(u6_mem_b0_b_96), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_120));
SDFFN u7_mem_reg_b2_b_b14_b (.CK(clk_i), .D(n_9014), .Q(u7_mem_b2_b_42), .SO(u7_mem_b2_b_42), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_96));
SDFFN u7_mem_reg_b2_b_b10_b (.CK(clk_i), .D(n_9019), .Q(u7_mem_b2_b_38), .SO(u7_mem_b2_b_38), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_42));
SDFFN u8_mem_reg_b2_b_b6_b (.CK(clk_i), .D(n_8473), .Q(u8_mem_b2_b_34), .SO(u8_mem_b2_b_34), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_38));
SDFFN u6_mem_reg_b0_b_b28_b (.CK(clk_i), .D(n_8763), .Q(u6_mem_b0_b_118), .SO(u6_mem_b0_b_118), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_34));
SDFFN u7_mem_reg_b1_b_b7_b (.CK(clk_i), .D(n_9025), .Q(u7_mem_b1_b_66), .SO(u7_mem_b1_b_66), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_118));
SDFFN u6_mem_reg_b3_b_b8_b (.CK(clk_i), .D(n_9074), .Q(u6_mem_b3_b_129), .SO(u6_mem_b3_b_129), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_66));
SDFFNSRN u13_crac_dout_r_reg_b3_b (.CK(clk_i), .D(n_8641), .Q(crac_out_848), .SO(crac_out_848), .SE(scan_enable), .SI(u6_mem_b3_b_129));
SDFFNSRN u13_crac_dout_r_reg_b9_b (.CK(clk_i), .D(n_8636), .Q(crac_out_854), .SO(crac_out_854), .SE(scan_enable), .SI(crac_out_848));
SDFFN u7_mem_reg_b1_b_b3_b (.CK(clk_i), .D(n_9030), .Q(u7_mem_b1_b_62), .SO(u7_mem_b1_b_62), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_out_854));
SDFFN u13_icc_r_reg_b22_b (.CK(clk_i), .D(n_8592), .Q(ic2_cfg_1049), .SO(ic2_cfg_1049), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_62));
SDFFNSRN u13_crac_dout_r_reg_b14_b (.CK(clk_i), .D(n_8649), .Q(crac_out_859), .SO(crac_out_859), .SE(scan_enable), .SI(ic2_cfg_1049));
SDFFN u13_occ0_r_reg_b2_b (.CK(clk_i), .D(n_8535), .Q(oc0_cfg_965), .SO(oc0_cfg_965), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_out_859));
SDFFN u13_occ0_r_reg_b4_b (.CK(clk_i), .D(n_8529), .Q(n_8528), .SO(n_8528), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc0_cfg_965));
SDFFN u13_intm_r_reg_b7_b (.CK(clk_i), .D(n_8489), .Q(u13_intm_r_b7_b), .SO(u13_intm_r_b7_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(n_8528));
SDFFN u13_intm_r_reg_b22_b (.CK(clk_i), .D(n_8506), .Q(u13_intm_r_b22_b), .SO(u13_intm_r_b22_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b7_b));
SDFFN u13_icc_r_reg_b11_b (.CK(clk_i), .D(n_8620), .Q(ic1_cfg_1036), .SO(ic1_cfg_1036), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b22_b));
SDFFN u7_mem_reg_b1_b_b29_b (.CK(clk_i), .D(n_9037), .Q(u7_mem_b1_b_88), .SO(u7_mem_b1_b_88), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic1_cfg_1036));
SDFFN u6_mem_reg_b0_b_b23_b (.CK(clk_i), .D(n_8767), .Q(u6_mem_b0_b_113), .SO(u6_mem_b0_b_113), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_88));
SDFFN u13_icc_r_reg_b15_b (.CK(clk_i), .D(n_8610), .Q(ic1_cfg_1040), .SO(ic1_cfg_1040), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_113));
SDFFN u13_icc_r_reg_b19_b (.CK(clk_i), .D(n_8601), .Q(ic2_cfg_1046), .SO(ic2_cfg_1046), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic1_cfg_1040));
SDFFN u13_crac_r_reg_b0_b (.CK(clk_i), .D(n_8635), .Q(crac_out_861), .SO(crac_out_861), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic2_cfg_1046));
SDFFN u13_crac_r_reg_b1_b (.CK(clk_i), .D(n_8633), .Q(crac_out_862), .SO(crac_out_862), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_out_861));
SDFFN u13_crac_r_reg_b3_b (.CK(clk_i), .D(n_8631), .Q(crac_out_864), .SO(crac_out_864), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_out_862));
SDFFN u13_crac_r_reg_b4_b (.CK(clk_i), .D(n_8630), .Q(crac_out_865), .SO(crac_out_865), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_out_864));
SDFFN u13_crac_r_reg_b5_b (.CK(clk_i), .D(n_8628), .Q(crac_out_866), .SO(crac_out_866), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_out_865));
SDFFN u13_crac_r_reg_b7_b (.CK(clk_i), .D(n_8626), .Q(crac_out_876), .SO(crac_out_876), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_out_866));
SDFFN u13_icc_r_reg_b0_b (.CK(clk_i), .D(n_8624), .Q(ic0_cfg), .SO(ic0_cfg), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_out_876));
SDFFN u13_icc_r_reg_b10_b (.CK(clk_i), .D(n_8622), .Q(ic1_cfg_1035), .SO(ic1_cfg_1035), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic0_cfg));
SDFFN u13_icc_r_reg_b12_b (.CK(clk_i), .D(n_8618), .Q(n_4736), .SO(n_4736), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic1_cfg_1035));
SDFFN u13_icc_r_reg_b13_b (.CK(clk_i), .D(n_8616), .Q(n_4734), .SO(n_4734), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(n_4736));
SDFFN u13_icc_r_reg_b14_b (.CK(clk_i), .D(n_8613), .Q(ic1_cfg_1039), .SO(ic1_cfg_1039), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(n_4734));
SDFFN u13_icc_r_reg_b16_b (.CK(clk_i), .D(n_8608), .Q(ic2_cfg), .SO(ic2_cfg), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic1_cfg_1039));
SDFFN u13_icc_r_reg_b17_b (.CK(clk_i), .D(n_8606), .Q(ic2_cfg_1044), .SO(ic2_cfg_1044), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic2_cfg));
SDFFN u13_icc_r_reg_b18_b (.CK(clk_i), .D(n_8604), .Q(ic2_cfg_1045), .SO(ic2_cfg_1045), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic2_cfg_1044));
SDFFN u13_icc_r_reg_b1_b (.CK(clk_i), .D(n_8599), .Q(ic0_cfg_1024), .SO(ic0_cfg_1024), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic2_cfg_1045));
SDFFN u13_icc_r_reg_b20_b (.CK(clk_i), .D(n_8597), .Q(n_5788), .SO(n_5788), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic0_cfg_1024));
SDFFN u13_icc_r_reg_b21_b (.CK(clk_i), .D(n_8594), .Q(n_5588), .SO(n_5588), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(n_5788));
SDFFN u13_icc_r_reg_b23_b (.CK(clk_i), .D(n_8589), .Q(ic2_cfg_1050), .SO(ic2_cfg_1050), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(n_5588));
SDFFN u13_icc_r_reg_b2_b (.CK(clk_i), .D(n_8588), .Q(ic0_cfg_1025), .SO(ic0_cfg_1025), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic2_cfg_1050));
SDFFN u13_icc_r_reg_b3_b (.CK(clk_i), .D(n_8586), .Q(ic0_cfg_1026), .SO(ic0_cfg_1026), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic0_cfg_1025));
SDFFN u13_icc_r_reg_b4_b (.CK(clk_i), .D(n_8584), .Q(n_4708), .SO(n_4708), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic0_cfg_1026));
SDFFN u13_icc_r_reg_b5_b (.CK(clk_i), .D(n_8581), .Q(n_4703), .SO(n_4703), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(n_4708));
SDFFN u13_icc_r_reg_b6_b (.CK(clk_i), .D(n_8579), .Q(ic0_cfg_1029), .SO(ic0_cfg_1029), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(n_4703));
SDFFN u13_icc_r_reg_b7_b (.CK(clk_i), .D(n_8577), .Q(ic0_cfg_1030), .SO(ic0_cfg_1030), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic0_cfg_1029));
SDFFN u13_icc_r_reg_b9_b (.CK(clk_i), .D(n_8573), .Q(ic1_cfg_1034), .SO(ic1_cfg_1034), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic0_cfg_1030));
SDFFN u13_occ0_r_reg_b0_b (.CK(clk_i), .D(n_8571), .Q(oc0_cfg), .SO(oc0_cfg), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic1_cfg_1034));
SDFFN u13_occ0_r_reg_b10_b (.CK(clk_i), .D(n_8570), .Q(oc1_cfg_975), .SO(oc1_cfg_975), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc0_cfg));
SDFFN u13_occ0_r_reg_b12_b (.CK(clk_i), .D(n_8568), .Q(n_8567), .SO(n_8567), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc1_cfg_975));
SDFFN u13_occ0_r_reg_b13_b (.CK(clk_i), .D(n_8566), .Q(n_8565), .SO(n_8565), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(n_8567));
SDFFN u13_occ0_r_reg_b14_b (.CK(clk_i), .D(n_8564), .Q(oc1_cfg_979), .SO(oc1_cfg_979), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(n_8565));
SDFFN u13_occ0_r_reg_b16_b (.CK(clk_i), .D(n_8562), .Q(oc2_cfg), .SO(oc2_cfg), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc1_cfg_979));
SDFFN u13_occ0_r_reg_b17_b (.CK(clk_i), .D(n_8560), .Q(oc2_cfg_984), .SO(oc2_cfg_984), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc2_cfg));
SDFFN u13_occ0_r_reg_b18_b (.CK(clk_i), .D(n_8558), .Q(oc2_cfg_985), .SO(oc2_cfg_985), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc2_cfg_984));
SDFFN u13_occ0_r_reg_b1_b (.CK(clk_i), .D(n_8555), .Q(oc0_cfg_964), .SO(oc0_cfg_964), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc2_cfg_985));
SDFFN u13_occ0_r_reg_b20_b (.CK(clk_i), .D(n_8554), .Q(oc2_cfg_987), .SO(oc2_cfg_987), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc0_cfg_964));
SDFFN u13_occ0_r_reg_b21_b (.CK(clk_i), .D(n_8551), .Q(n_8550), .SO(n_8550), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc2_cfg_987));
SDFFN u13_occ0_r_reg_b23_b (.CK(clk_i), .D(n_8548), .Q(oc2_cfg_990), .SO(oc2_cfg_990), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(n_8550));
SDFFN u13_occ0_r_reg_b24_b (.CK(clk_i), .D(n_8546), .Q(oc3_cfg), .SO(oc3_cfg), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc2_cfg_990));
SDFFN u13_occ0_r_reg_b25_b (.CK(clk_i), .D(n_8545), .Q(oc3_cfg_994), .SO(oc3_cfg_994), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc3_cfg));
SDFFN u13_occ0_r_reg_b27_b (.CK(clk_i), .D(n_8542), .Q(oc3_cfg_996), .SO(oc3_cfg_996), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc3_cfg_994));
SDFFN u13_occ0_r_reg_b28_b (.CK(clk_i), .D(n_8540), .Q(oc3_cfg_997), .SO(oc3_cfg_997), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc3_cfg_996));
SDFFN u13_occ0_r_reg_b29_b (.CK(clk_i), .D(n_8537), .Q(n_8536), .SO(n_8536), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc3_cfg_997));
SDFFN u13_occ0_r_reg_b30_b (.CK(clk_i), .D(n_8534), .Q(oc3_cfg_999), .SO(oc3_cfg_999), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(n_8536));
SDFFN u13_occ0_r_reg_b31_b (.CK(clk_i), .D(n_8532), .Q(oc3_cfg_1000), .SO(oc3_cfg_1000), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc3_cfg_999));
SDFFN u13_occ0_r_reg_b3_b (.CK(clk_i), .D(n_8530), .Q(oc0_cfg_966), .SO(oc0_cfg_966), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc3_cfg_1000));
SDFFN u13_occ0_r_reg_b5_b (.CK(clk_i), .D(n_8527), .Q(n_8526), .SO(n_8526), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc0_cfg_966));
SDFFN u13_occ0_r_reg_b6_b (.CK(clk_i), .D(n_8525), .Q(oc0_cfg_969), .SO(oc0_cfg_969), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(n_8526));
SDFFN u13_occ0_r_reg_b7_b (.CK(clk_i), .D(n_8524), .Q(oc0_cfg_970), .SO(oc0_cfg_970), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc0_cfg_969));
SDFFN u13_occ0_r_reg_b9_b (.CK(clk_i), .D(n_8522), .Q(oc1_cfg_974), .SO(oc1_cfg_974), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc0_cfg_970));
SDFFN u13_intm_r_reg_b0_b (.CK(clk_i), .D(n_8521), .Q(u13_intm_r_b0_b), .SO(u13_intm_r_b0_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc1_cfg_974));
SDFFN u13_intm_r_reg_b10_b (.CK(clk_i), .D(n_8520), .Q(u13_intm_r_b10_b), .SO(u13_intm_r_b10_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b0_b));
SDFFN u13_intm_r_reg_b11_b (.CK(clk_i), .D(n_8518), .Q(u13_intm_r_b11_b), .SO(u13_intm_r_b11_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b10_b));
SDFFN u13_intm_r_reg_b12_b (.CK(clk_i), .D(n_8517), .Q(u13_intm_r_b12_b), .SO(u13_intm_r_b12_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b11_b));
SDFFN u13_intm_r_reg_b13_b (.CK(clk_i), .D(n_8516), .Q(u13_intm_r_b13_b), .SO(u13_intm_r_b13_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b12_b));
SDFFN u13_intm_r_reg_b14_b (.CK(clk_i), .D(n_8515), .Q(u13_intm_r_b14_b), .SO(u13_intm_r_b14_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b13_b));
SDFFN u13_intm_r_reg_b16_b (.CK(clk_i), .D(n_8513), .Q(u13_intm_r_b16_b), .SO(u13_intm_r_b16_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b14_b));
SDFFN u13_intm_r_reg_b17_b (.CK(clk_i), .D(n_8512), .Q(u13_intm_r_b17_b), .SO(u13_intm_r_b17_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b16_b));
SDFFN u13_intm_r_reg_b18_b (.CK(clk_i), .D(n_8511), .Q(u13_intm_r_b18_b), .SO(u13_intm_r_b18_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b17_b));
SDFFN u13_intm_r_reg_b19_b (.CK(clk_i), .D(n_8510), .Q(u13_intm_r_b19_b), .SO(u13_intm_r_b19_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b18_b));
SDFFN u13_intm_r_reg_b1_b (.CK(clk_i), .D(n_8509), .Q(u13_intm_r_b1_b), .SO(u13_intm_r_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b19_b));
SDFFN u13_intm_r_reg_b20_b (.CK(clk_i), .D(n_8508), .Q(u13_intm_r_b20_b), .SO(u13_intm_r_b20_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b1_b));
SDFFN u13_intm_r_reg_b21_b (.CK(clk_i), .D(n_8507), .Q(u13_intm_r_b21_b), .SO(u13_intm_r_b21_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b20_b));
SDFFN u13_intm_r_reg_b23_b (.CK(clk_i), .D(n_8505), .Q(u13_intm_r_b23_b), .SO(u13_intm_r_b23_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b21_b));
SDFFN u13_intm_r_reg_b24_b (.CK(clk_i), .D(n_8504), .Q(u13_intm_r_b24_b), .SO(u13_intm_r_b24_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b23_b));
SDFFN u13_intm_r_reg_b25_b (.CK(clk_i), .D(n_8502), .Q(u13_intm_r_b25_b), .SO(u13_intm_r_b25_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b24_b));
SDFFN u13_intm_r_reg_b27_b (.CK(clk_i), .D(n_8498), .Q(u13_intm_r_b27_b), .SO(u13_intm_r_b27_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b25_b));
SDFFN u13_intm_r_reg_b28_b (.CK(clk_i), .D(n_8496), .Q(u13_intm_r_b28_b), .SO(u13_intm_r_b28_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b27_b));
SDFFN u13_intm_r_reg_b2_b (.CK(clk_i), .D(n_8494), .Q(u13_intm_r_b2_b), .SO(u13_intm_r_b2_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b28_b));
SDFFN u13_intm_r_reg_b5_b (.CK(clk_i), .D(n_8491), .Q(u13_intm_r_b5_b), .SO(u13_intm_r_b5_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b2_b));
SDFFN u13_intm_r_reg_b6_b (.CK(clk_i), .D(n_8490), .Q(u13_intm_r_b6_b), .SO(u13_intm_r_b6_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b5_b));
SDFFN u13_intm_r_reg_b9_b (.CK(clk_i), .D(n_8487), .Q(u13_intm_r_b9_b), .SO(u13_intm_r_b9_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b6_b));
SDFFN u13_intm_r_reg_b4_b (.CK(clk_i), .D(n_8492), .Q(u13_intm_r_b4_b), .SO(u13_intm_r_b4_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b9_b));
SDFFN u13_intm_r_reg_b15_b (.CK(clk_i), .D(n_8514), .Q(u13_intm_r_b15_b), .SO(u13_intm_r_b15_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b4_b));
SDFFNSRN u13_crac_dout_r_reg_b0_b (.CK(clk_i), .D(n_8655), .Q(crac_out), .SO(crac_out), .SE(scan_enable), .SI(u13_intm_r_b15_b));
SDFFNSRN u13_crac_dout_r_reg_b10_b (.CK(clk_i), .D(n_8654), .Q(crac_out_855), .SO(crac_out_855), .SE(scan_enable), .SI(crac_out));
SDFFNSRN u13_crac_dout_r_reg_b11_b (.CK(clk_i), .D(n_8653), .Q(crac_out_856), .SO(crac_out_856), .SE(scan_enable), .SI(crac_out_855));
SDFFNSRN u13_crac_dout_r_reg_b12_b (.CK(clk_i), .D(n_8652), .Q(crac_out_857), .SO(crac_out_857), .SE(scan_enable), .SI(crac_out_856));
SDFFNSRN u13_crac_dout_r_reg_b13_b (.CK(clk_i), .D(n_8651), .Q(crac_out_858), .SO(crac_out_858), .SE(scan_enable), .SI(crac_out_857));
SDFFNSRN u13_crac_dout_r_reg_b15_b (.CK(clk_i), .D(n_8648), .Q(crac_out_860), .SO(crac_out_860), .SE(scan_enable), .SI(crac_out_858));
SDFFNSRN u13_crac_dout_r_reg_b1_b (.CK(clk_i), .D(n_8646), .Q(crac_out_846), .SO(crac_out_846), .SE(scan_enable), .SI(crac_out_860));
SDFFNSRN u13_crac_dout_r_reg_b2_b (.CK(clk_i), .D(n_8644), .Q(crac_out_847), .SO(crac_out_847), .SE(scan_enable), .SI(crac_out_846));
SDFFNSRN u13_crac_dout_r_reg_b4_b (.CK(clk_i), .D(n_8642), .Q(crac_out_849), .SO(crac_out_849), .SE(scan_enable), .SI(crac_out_847));
SDFFNSRN u13_crac_dout_r_reg_b5_b (.CK(clk_i), .D(n_8640), .Q(crac_out_850), .SO(crac_out_850), .SE(scan_enable), .SI(crac_out_849));
SDFFNSRN u13_crac_dout_r_reg_b6_b (.CK(clk_i), .D(n_8639), .Q(crac_out_851), .SO(crac_out_851), .SE(scan_enable), .SI(crac_out_850));
SDFFNSRN u13_crac_dout_r_reg_b8_b (.CK(clk_i), .D(n_8637), .Q(crac_out_853), .SO(crac_out_853), .SE(scan_enable), .SI(crac_out_851));
SDFFN u8_mem_reg_b2_b_b4_b (.CK(clk_i), .D(n_8845), .Q(u8_mem_b2_b_32), .SO(u8_mem_b2_b_32), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_out_853));
SDFFN u3_mem_reg_b1_b_b28_b (.CK(clk_i), .D(n_8846), .Q(u3_mem_b1_b_87), .SO(u3_mem_b1_b_87), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_32));
SDFFN u8_mem_reg_b2_b_b5_b (.CK(clk_i), .D(n_8475), .Q(u8_mem_b2_b_33), .SO(u8_mem_b2_b_33), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_87));
SDFFN u3_mem_reg_b1_b_b29_b (.CK(clk_i), .D(n_8474), .Q(u3_mem_b1_b_88), .SO(u3_mem_b1_b_88), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_33));
SDFFN u8_mem_reg_b2_b_b7_b (.CK(clk_i), .D(n_8472), .Q(u8_mem_b2_b_35), .SO(u8_mem_b2_b_35), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_88));
SDFFN u8_mem_reg_b2_b_b8_b (.CK(clk_i), .D(n_8470), .Q(u8_mem_b2_b_36), .SO(u8_mem_b2_b_36), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_35));
SDFFN u8_mem_reg_b2_b_b9_b (.CK(clk_i), .D(n_8469), .Q(u8_mem_b2_b_37), .SO(u8_mem_b2_b_37), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_36));
SDFFN u8_mem_reg_b3_b_b0_b (.CK(clk_i), .D(n_8467), .Q(u8_mem_b3_b), .SO(u8_mem_b3_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_37));
SDFFN u3_mem_reg_b1_b_b30_b (.CK(clk_i), .D(n_8408), .Q(u3_mem_b1_b_89), .SO(u3_mem_b1_b_89), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b));
SDFFN u8_mem_reg_b3_b_b11_b (.CK(clk_i), .D(n_8903), .Q(u8_mem_b3_b_132), .SO(u8_mem_b3_b_132), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_89));
SDFFN u3_mem_reg_b1_b_b31_b (.CK(clk_i), .D(n_8463), .Q(u3_mem_b1_b_90), .SO(u3_mem_b1_b_90), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_132));
SDFFN u8_mem_reg_b3_b_b12_b (.CK(clk_i), .D(n_8462), .Q(u8_mem_b3_b_133), .SO(u8_mem_b3_b_133), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_90));
SDFFN u8_mem_reg_b3_b_b13_b (.CK(clk_i), .D(n_8459), .Q(u8_mem_b3_b_134), .SO(u8_mem_b3_b_134), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_133));
SDFFN u3_mem_reg_b1_b_b4_b (.CK(clk_i), .D(n_8455), .Q(u3_mem_b1_b_63), .SO(u3_mem_b1_b_63), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_134));
SDFFN u8_mem_reg_b3_b_b14_b (.CK(clk_i), .D(n_8458), .Q(u8_mem_b3_b_135), .SO(u8_mem_b3_b_135), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_63));
SDFFN u8_mem_reg_b3_b_b16_b (.CK(clk_i), .D(n_8454), .Q(u8_mem_b3_b_137), .SO(u8_mem_b3_b_137), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_135));
SDFFN u8_mem_reg_b3_b_b17_b (.CK(clk_i), .D(n_8450), .Q(u8_mem_b3_b_138), .SO(u8_mem_b3_b_138), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_137));
SDFFN u3_mem_reg_b1_b_b5_b (.CK(clk_i), .D(n_8452), .Q(u3_mem_b1_b_64), .SO(u3_mem_b1_b_64), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_138));
SDFFN u8_mem_reg_b3_b_b19_b (.CK(clk_i), .D(n_8468), .Q(u8_mem_b3_b_140), .SO(u8_mem_b3_b_140), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_64));
SDFFN u3_mem_reg_b1_b_b6_b (.CK(clk_i), .D(n_8447), .Q(u3_mem_b1_b_65), .SO(u3_mem_b1_b_65), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_140));
SDFFN u8_mem_reg_b3_b_b1_b (.CK(clk_i), .D(n_8446), .Q(u8_mem_b3_b_122), .SO(u8_mem_b3_b_122), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_65));
SDFFN u3_mem_reg_b1_b_b7_b (.CK(clk_i), .D(n_8445), .Q(u3_mem_b1_b_66), .SO(u3_mem_b1_b_66), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_122));
SDFFN u8_mem_reg_b3_b_b20_b (.CK(clk_i), .D(n_8443), .Q(u8_mem_b3_b_141), .SO(u8_mem_b3_b_141), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_66));
SDFFN u8_mem_reg_b3_b_b21_b (.CK(clk_i), .D(n_8442), .Q(u8_mem_b3_b_142), .SO(u8_mem_b3_b_142), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_141));
SDFFN u3_mem_reg_b1_b_b8_b (.CK(clk_i), .D(n_8441), .Q(u3_mem_b1_b_67), .SO(u3_mem_b1_b_67), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_142));
SDFFN u8_mem_reg_b3_b_b23_b (.CK(clk_i), .D(n_8437), .Q(u8_mem_b3_b_144), .SO(u8_mem_b3_b_144), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_67));
SDFFN u8_mem_reg_b3_b_b24_b (.CK(clk_i), .D(n_8435), .Q(u8_mem_b3_b_145), .SO(u8_mem_b3_b_145), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_144));
SDFFN u3_mem_reg_b1_b_b9_b (.CK(clk_i), .D(n_8436), .Q(u3_mem_b1_b_68), .SO(u3_mem_b1_b_68), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_145));
SDFFN u8_mem_reg_b3_b_b26_b (.CK(clk_i), .D(n_8350), .Q(u8_mem_b3_b_147), .SO(u8_mem_b3_b_147), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_68));
SDFFN u3_mem_reg_b2_b_b0_b (.CK(clk_i), .D(n_8432), .Q(u3_mem_b2_b), .SO(u3_mem_b2_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_147));
SDFFN u8_mem_reg_b3_b_b27_b (.CK(clk_i), .D(n_8431), .Q(u8_mem_b3_b_148), .SO(u8_mem_b3_b_148), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b));
SDFFN u3_mem_reg_b2_b_b10_b (.CK(clk_i), .D(n_8430), .Q(u3_mem_b2_b_38), .SO(u3_mem_b2_b_38), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_148));
SDFFN u8_mem_reg_b3_b_b29_b (.CK(clk_i), .D(n_8428), .Q(u8_mem_b3_b_150), .SO(u8_mem_b3_b_150), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_38));
SDFFN u8_mem_reg_b3_b_b2_b (.CK(clk_i), .D(n_8426), .Q(u8_mem_b3_b_123), .SO(u8_mem_b3_b_123), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_150));
SDFFN u8_mem_reg_b3_b_b30_b (.CK(clk_i), .D(n_8425), .Q(u8_mem_b3_b_151), .SO(u8_mem_b3_b_151), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_123));
SDFFN u8_mem_reg_b3_b_b31_b (.CK(clk_i), .D(n_9193), .Q(u8_mem_b3_b_152), .SO(u8_mem_b3_b_152), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_151));
SDFFN u3_mem_reg_b2_b_b12_b (.CK(clk_i), .D(n_8424), .Q(u3_mem_b2_b_40), .SO(u3_mem_b2_b_40), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_152));
SDFFN u8_mem_reg_b3_b_b4_b (.CK(clk_i), .D(n_9070), .Q(u8_mem_b3_b_125), .SO(u8_mem_b3_b_125), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_40));
SDFFN u3_mem_reg_b2_b_b13_b (.CK(clk_i), .D(n_8421), .Q(u3_mem_b2_b_41), .SO(u3_mem_b2_b_41), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_125));
SDFFN u8_mem_reg_b3_b_b5_b (.CK(clk_i), .D(n_8420), .Q(u8_mem_b3_b_126), .SO(u8_mem_b3_b_126), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_41));
SDFFN u3_mem_reg_b2_b_b14_b (.CK(clk_i), .D(n_9318), .Q(u3_mem_b2_b_42), .SO(u3_mem_b2_b_42), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_126));
SDFFN u8_mem_reg_b3_b_b7_b (.CK(clk_i), .D(n_8419), .Q(u8_mem_b3_b_128), .SO(u8_mem_b3_b_128), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_42));
SDFFN u3_mem_reg_b2_b_b15_b (.CK(clk_i), .D(n_8418), .Q(u3_mem_b2_b_43), .SO(u3_mem_b2_b_43), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_128));
SDFFN u8_mem_reg_b3_b_b9_b (.CK(clk_i), .D(n_8416), .Q(u8_mem_b3_b_130), .SO(u8_mem_b3_b_130), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_43));
SDFFN u3_mem_reg_b2_b_b16_b (.CK(clk_i), .D(n_8415), .Q(u3_mem_b2_b_44), .SO(u3_mem_b2_b_44), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b3_b_130));
SDFFN u3_mem_reg_b2_b_b17_b (.CK(clk_i), .D(n_8943), .Q(u3_mem_b2_b_45), .SO(u3_mem_b2_b_45), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_44));
SDFFN u3_mem_reg_b2_b_b19_b (.CK(clk_i), .D(n_8411), .Q(u3_mem_b2_b_47), .SO(u3_mem_b2_b_47), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_45));
SDFFN u3_mem_reg_b2_b_b1_b (.CK(clk_i), .D(n_8410), .Q(u3_mem_b2_b_29), .SO(u3_mem_b2_b_29), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_47));
SDFFN u3_mem_reg_b2_b_b21_b (.CK(clk_i), .D(n_8407), .Q(u3_mem_b2_b_49), .SO(u3_mem_b2_b_49), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_29));
SDFFN u3_mem_reg_b2_b_b23_b (.CK(clk_i), .D(n_8346), .Q(u3_mem_b2_b_51), .SO(u3_mem_b2_b_51), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_49));
SDFFN u3_mem_reg_b2_b_b24_b (.CK(clk_i), .D(n_8405), .Q(u3_mem_b2_b_52), .SO(u3_mem_b2_b_52), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_51));
SDFFN u3_mem_reg_b2_b_b25_b (.CK(clk_i), .D(n_9071), .Q(u3_mem_b2_b_53), .SO(u3_mem_b2_b_53), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_52));
SDFFN u3_mem_reg_b2_b_b27_b (.CK(clk_i), .D(n_8403), .Q(u3_mem_b2_b_55), .SO(u3_mem_b2_b_55), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_53));
SDFFN u3_mem_reg_b2_b_b28_b (.CK(clk_i), .D(n_8402), .Q(u3_mem_b2_b_56), .SO(u3_mem_b2_b_56), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_55));
SDFFN u3_mem_reg_b2_b_b29_b (.CK(clk_i), .D(n_8401), .Q(u3_mem_b2_b_57), .SO(u3_mem_b2_b_57), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_56));
SDFFN u3_mem_reg_b2_b_b30_b (.CK(clk_i), .D(n_8399), .Q(u3_mem_b2_b_58), .SO(u3_mem_b2_b_58), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_57));
SDFFN u3_mem_reg_b2_b_b31_b (.CK(clk_i), .D(n_8398), .Q(u3_mem_b2_b_59), .SO(u3_mem_b2_b_59), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_58));
SDFFN u3_mem_reg_b2_b_b3_b (.CK(clk_i), .D(n_8397), .Q(u3_mem_b2_b_31), .SO(u3_mem_b2_b_31), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_59));
SDFFN u3_mem_reg_b2_b_b4_b (.CK(clk_i), .D(n_8396), .Q(u3_mem_b2_b_32), .SO(u3_mem_b2_b_32), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_31));
SDFFN u3_mem_reg_b2_b_b5_b (.CK(clk_i), .D(n_8395), .Q(u3_mem_b2_b_33), .SO(u3_mem_b2_b_33), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_32));
SDFFN u3_mem_reg_b2_b_b6_b (.CK(clk_i), .D(n_8394), .Q(u3_mem_b2_b_34), .SO(u3_mem_b2_b_34), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_33));
SDFFN u3_mem_reg_b2_b_b7_b (.CK(clk_i), .D(n_8392), .Q(u3_mem_b2_b_35), .SO(u3_mem_b2_b_35), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_34));
SDFFN u3_mem_reg_b2_b_b9_b (.CK(clk_i), .D(n_8390), .Q(u3_mem_b2_b_37), .SO(u3_mem_b2_b_37), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_35));
SDFFN u3_mem_reg_b3_b_b0_b (.CK(clk_i), .D(n_8389), .Q(u3_mem_b3_b), .SO(u3_mem_b3_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_37));
SDFFN u3_mem_reg_b3_b_b10_b (.CK(clk_i), .D(n_8388), .Q(u3_mem_b3_b_131), .SO(u3_mem_b3_b_131), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b));
SDFFN u3_mem_reg_b3_b_b12_b (.CK(clk_i), .D(n_8385), .Q(u3_mem_b3_b_133), .SO(u3_mem_b3_b_133), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_131));
SDFFN u3_mem_reg_b3_b_b13_b (.CK(clk_i), .D(n_8384), .Q(u3_mem_b3_b_134), .SO(u3_mem_b3_b_134), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_133));
SDFFN u3_mem_reg_b3_b_b14_b (.CK(clk_i), .D(n_8382), .Q(u3_mem_b3_b_135), .SO(u3_mem_b3_b_135), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_134));
SDFFN u3_mem_reg_b3_b_b16_b (.CK(clk_i), .D(n_8379), .Q(u3_mem_b3_b_137), .SO(u3_mem_b3_b_137), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_135));
SDFFN u3_mem_reg_b3_b_b17_b (.CK(clk_i), .D(n_8378), .Q(u3_mem_b3_b_138), .SO(u3_mem_b3_b_138), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_137));
SDFFN u3_mem_reg_b3_b_b18_b (.CK(clk_i), .D(n_8377), .Q(u3_mem_b3_b_139), .SO(u3_mem_b3_b_139), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_138));
SDFFN u3_mem_reg_b3_b_b1_b (.CK(clk_i), .D(n_8374), .Q(u3_mem_b3_b_122), .SO(u3_mem_b3_b_122), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_139));
SDFFN u3_mem_reg_b3_b_b20_b (.CK(clk_i), .D(n_9023), .Q(u3_mem_b3_b_141), .SO(u3_mem_b3_b_141), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_122));
SDFFN u3_mem_reg_b3_b_b21_b (.CK(clk_i), .D(n_8373), .Q(u3_mem_b3_b_142), .SO(u3_mem_b3_b_142), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_141));
SDFFN u3_mem_reg_b3_b_b23_b (.CK(clk_i), .D(n_8370), .Q(u3_mem_b3_b_144), .SO(u3_mem_b3_b_144), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_142));
SDFFN u3_mem_reg_b3_b_b24_b (.CK(clk_i), .D(n_8368), .Q(u3_mem_b3_b_145), .SO(u3_mem_b3_b_145), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_144));
SDFFN u3_mem_reg_b3_b_b26_b (.CK(clk_i), .D(n_8367), .Q(u3_mem_b3_b_147), .SO(u3_mem_b3_b_147), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_145));
SDFFN u3_mem_reg_b3_b_b28_b (.CK(clk_i), .D(n_8364), .Q(u3_mem_b3_b_149), .SO(u3_mem_b3_b_149), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_147));
SDFFN u3_mem_reg_b3_b_b29_b (.CK(clk_i), .D(n_8363), .Q(u3_mem_b3_b_150), .SO(u3_mem_b3_b_150), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_149));
SDFFN u3_mem_reg_b3_b_b2_b (.CK(clk_i), .D(n_8362), .Q(u3_mem_b3_b_123), .SO(u3_mem_b3_b_123), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_150));
SDFFN u3_mem_reg_b3_b_b31_b (.CK(clk_i), .D(n_8360), .Q(u3_mem_b3_b_152), .SO(u3_mem_b3_b_152), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_123));
SDFFN u3_mem_reg_b3_b_b4_b (.CK(clk_i), .D(n_8359), .Q(u3_mem_b3_b_125), .SO(u3_mem_b3_b_125), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_152));
SDFFN u3_mem_reg_b3_b_b5_b (.CK(clk_i), .D(n_8358), .Q(u3_mem_b3_b_126), .SO(u3_mem_b3_b_126), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_125));
SDFFN u3_mem_reg_b3_b_b7_b (.CK(clk_i), .D(n_8354), .Q(u3_mem_b3_b_128), .SO(u3_mem_b3_b_128), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_126));
SDFFN u3_mem_reg_b3_b_b9_b (.CK(clk_i), .D(n_8352), .Q(u3_mem_b3_b_130), .SO(u3_mem_b3_b_130), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_128));
SDFFN u3_mem_reg_b3_b_b25_b (.CK(clk_i), .D(n_8348), .Q(u3_mem_b3_b_146), .SO(u3_mem_b3_b_146), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_130));
SDFFN u4_mem_reg_b1_b_b0_b (.CK(clk_i), .D(n_8345), .Q(u4_mem_b1_b), .SO(u4_mem_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_146));
SDFFN u4_mem_reg_b1_b_b10_b (.CK(clk_i), .D(n_8344), .Q(u4_mem_b1_b_69), .SO(u4_mem_b1_b_69), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b));
SDFFN u4_mem_reg_b1_b_b11_b (.CK(clk_i), .D(n_8343), .Q(u4_mem_b1_b_70), .SO(u4_mem_b1_b_70), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_69));
SDFFN u4_mem_reg_b1_b_b13_b (.CK(clk_i), .D(n_8341), .Q(u4_mem_b1_b_72), .SO(u4_mem_b1_b_72), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_70));
SDFFN u4_mem_reg_b1_b_b14_b (.CK(clk_i), .D(n_8340), .Q(u4_mem_b1_b_73), .SO(u4_mem_b1_b_73), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_72));
SDFFN u4_mem_reg_b1_b_b15_b (.CK(clk_i), .D(n_8338), .Q(u4_mem_b1_b_74), .SO(u4_mem_b1_b_74), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_73));
SDFFN u4_mem_reg_b1_b_b17_b (.CK(clk_i), .D(n_8334), .Q(u4_mem_b1_b_76), .SO(u4_mem_b1_b_76), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_74));
SDFFN u4_mem_reg_b1_b_b18_b (.CK(clk_i), .D(n_8332), .Q(u4_mem_b1_b_77), .SO(u4_mem_b1_b_77), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_76));
SDFFN u4_mem_reg_b1_b_b19_b (.CK(clk_i), .D(n_8330), .Q(u4_mem_b1_b_78), .SO(u4_mem_b1_b_78), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_77));
SDFFN u4_mem_reg_b1_b_b1_b (.CK(clk_i), .D(n_8329), .Q(u4_mem_b1_b_60), .SO(u4_mem_b1_b_60), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_78));
SDFFN u4_mem_reg_b1_b_b20_b (.CK(clk_i), .D(n_8328), .Q(u4_mem_b1_b_79), .SO(u4_mem_b1_b_79), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_60));
SDFFN u4_mem_reg_b1_b_b21_b (.CK(clk_i), .D(n_8327), .Q(u4_mem_b1_b_80), .SO(u4_mem_b1_b_80), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_79));
SDFFN u4_mem_reg_b1_b_b22_b (.CK(clk_i), .D(n_8326), .Q(u4_mem_b1_b_81), .SO(u4_mem_b1_b_81), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_80));
SDFFN u4_mem_reg_b1_b_b24_b (.CK(clk_i), .D(n_8324), .Q(u4_mem_b1_b_83), .SO(u4_mem_b1_b_83), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_81));
SDFFN u4_mem_reg_b1_b_b25_b (.CK(clk_i), .D(n_8322), .Q(u4_mem_b1_b_84), .SO(u4_mem_b1_b_84), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_83));
SDFFN u4_mem_reg_b1_b_b26_b (.CK(clk_i), .D(n_8321), .Q(u4_mem_b1_b_85), .SO(u4_mem_b1_b_85), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_84));
SDFFN u4_mem_reg_b1_b_b28_b (.CK(clk_i), .D(n_8319), .Q(u4_mem_b1_b_87), .SO(u4_mem_b1_b_87), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_85));
SDFFN u4_mem_reg_b1_b_b29_b (.CK(clk_i), .D(n_8317), .Q(u4_mem_b1_b_88), .SO(u4_mem_b1_b_88), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_87));
SDFFN u4_mem_reg_b1_b_b2_b (.CK(clk_i), .D(n_8315), .Q(u4_mem_b1_b_61), .SO(u4_mem_b1_b_61), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_88));
SDFFN u4_mem_reg_b1_b_b31_b (.CK(clk_i), .D(n_8311), .Q(u4_mem_b1_b_90), .SO(u4_mem_b1_b_90), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_61));
SDFFN u4_mem_reg_b1_b_b3_b (.CK(clk_i), .D(n_8310), .Q(u4_mem_b1_b_62), .SO(u4_mem_b1_b_62), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_90));
SDFFN u4_mem_reg_b1_b_b4_b (.CK(clk_i), .D(n_8309), .Q(u4_mem_b1_b_63), .SO(u4_mem_b1_b_63), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_62));
SDFFN u4_mem_reg_b1_b_b6_b (.CK(clk_i), .D(n_8306), .Q(u4_mem_b1_b_65), .SO(u4_mem_b1_b_65), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_63));
SDFFN u4_mem_reg_b1_b_b7_b (.CK(clk_i), .D(n_8305), .Q(u4_mem_b1_b_66), .SO(u4_mem_b1_b_66), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_65));
SDFFN u4_mem_reg_b1_b_b8_b (.CK(clk_i), .D(n_8304), .Q(u4_mem_b1_b_67), .SO(u4_mem_b1_b_67), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_66));
SDFFN u4_mem_reg_b2_b_b0_b (.CK(clk_i), .D(n_8302), .Q(u4_mem_b2_b), .SO(u4_mem_b2_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b1_b_67));
SDFFN u4_mem_reg_b2_b_b10_b (.CK(clk_i), .D(n_8301), .Q(u4_mem_b2_b_38), .SO(u4_mem_b2_b_38), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b));
SDFFN u4_mem_reg_b2_b_b11_b (.CK(clk_i), .D(n_8300), .Q(u4_mem_b2_b_39), .SO(u4_mem_b2_b_39), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_38));
SDFFN u4_mem_reg_b2_b_b13_b (.CK(clk_i), .D(n_8297), .Q(u4_mem_b2_b_41), .SO(u4_mem_b2_b_41), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_39));
SDFFN u4_mem_reg_b2_b_b14_b (.CK(clk_i), .D(n_8296), .Q(u4_mem_b2_b_42), .SO(u4_mem_b2_b_42), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_41));
SDFFN u4_mem_reg_b2_b_b15_b (.CK(clk_i), .D(n_8295), .Q(u4_mem_b2_b_43), .SO(u4_mem_b2_b_43), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_42));
SDFFN u4_mem_reg_b2_b_b17_b (.CK(clk_i), .D(n_8293), .Q(u4_mem_b2_b_45), .SO(u4_mem_b2_b_45), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_43));
SDFFN u4_mem_reg_b2_b_b18_b (.CK(clk_i), .D(n_8291), .Q(u4_mem_b2_b_46), .SO(u4_mem_b2_b_46), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_45));
SDFFN u4_mem_reg_b2_b_b19_b (.CK(clk_i), .D(n_8290), .Q(u4_mem_b2_b_47), .SO(u4_mem_b2_b_47), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_46));
SDFFN u4_mem_reg_b2_b_b1_b (.CK(clk_i), .D(n_8289), .Q(u4_mem_b2_b_29), .SO(u4_mem_b2_b_29), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_47));
SDFFN u4_mem_reg_b2_b_b20_b (.CK(clk_i), .D(n_8287), .Q(u4_mem_b2_b_48), .SO(u4_mem_b2_b_48), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_29));
SDFFN u4_mem_reg_b2_b_b21_b (.CK(clk_i), .D(n_8286), .Q(u4_mem_b2_b_49), .SO(u4_mem_b2_b_49), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_48));
SDFFN u4_mem_reg_b2_b_b22_b (.CK(clk_i), .D(n_8285), .Q(u4_mem_b2_b_50), .SO(u4_mem_b2_b_50), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_49));
SDFFN u4_mem_reg_b2_b_b24_b (.CK(clk_i), .D(n_8283), .Q(u4_mem_b2_b_52), .SO(u4_mem_b2_b_52), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_50));
SDFFN u4_mem_reg_b2_b_b25_b (.CK(clk_i), .D(n_8282), .Q(u4_mem_b2_b_53), .SO(u4_mem_b2_b_53), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_52));
SDFFN u4_mem_reg_b2_b_b26_b (.CK(clk_i), .D(n_8281), .Q(u4_mem_b2_b_54), .SO(u4_mem_b2_b_54), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_53));
SDFFN u4_mem_reg_b2_b_b28_b (.CK(clk_i), .D(n_8278), .Q(u4_mem_b2_b_56), .SO(u4_mem_b2_b_56), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_54));
SDFFN u4_mem_reg_b2_b_b29_b (.CK(clk_i), .D(n_8277), .Q(u4_mem_b2_b_57), .SO(u4_mem_b2_b_57), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_56));
SDFFN u4_mem_reg_b2_b_b2_b (.CK(clk_i), .D(n_8275), .Q(u4_mem_b2_b_30), .SO(u4_mem_b2_b_30), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_57));
SDFFN u4_mem_reg_b2_b_b31_b (.CK(clk_i), .D(n_8273), .Q(u4_mem_b2_b_59), .SO(u4_mem_b2_b_59), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_30));
SDFFN u4_mem_reg_b2_b_b3_b (.CK(clk_i), .D(n_8272), .Q(u4_mem_b2_b_31), .SO(u4_mem_b2_b_31), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_59));
SDFFN u4_mem_reg_b2_b_b4_b (.CK(clk_i), .D(n_8271), .Q(u4_mem_b2_b_32), .SO(u4_mem_b2_b_32), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_31));
SDFFN u4_mem_reg_b2_b_b6_b (.CK(clk_i), .D(n_8269), .Q(u4_mem_b2_b_34), .SO(u4_mem_b2_b_34), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_32));
SDFFN u4_mem_reg_b2_b_b7_b (.CK(clk_i), .D(n_8268), .Q(u4_mem_b2_b_35), .SO(u4_mem_b2_b_35), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_34));
SDFFN u4_mem_reg_b2_b_b8_b (.CK(clk_i), .D(n_8267), .Q(u4_mem_b2_b_36), .SO(u4_mem_b2_b_36), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_35));
SDFFN u4_mem_reg_b3_b_b0_b (.CK(clk_i), .D(n_8265), .Q(u4_mem_b3_b), .SO(u4_mem_b3_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b2_b_36));
SDFFN u4_mem_reg_b3_b_b10_b (.CK(clk_i), .D(n_8264), .Q(u4_mem_b3_b_131), .SO(u4_mem_b3_b_131), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b));
SDFFN u4_mem_reg_b3_b_b11_b (.CK(clk_i), .D(n_8262), .Q(u4_mem_b3_b_132), .SO(u4_mem_b3_b_132), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_131));
SDFFN u4_mem_reg_b3_b_b13_b (.CK(clk_i), .D(n_8260), .Q(u4_mem_b3_b_134), .SO(u4_mem_b3_b_134), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_132));
SDFFN u4_mem_reg_b3_b_b14_b (.CK(clk_i), .D(n_8259), .Q(u4_mem_b3_b_135), .SO(u4_mem_b3_b_135), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_134));
SDFFN u4_mem_reg_b3_b_b15_b (.CK(clk_i), .D(n_9351), .Q(u4_mem_b3_b_136), .SO(u4_mem_b3_b_136), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_135));
SDFFN u4_mem_reg_b3_b_b17_b (.CK(clk_i), .D(n_9348), .Q(u4_mem_b3_b_138), .SO(u4_mem_b3_b_138), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_136));
SDFFN u4_mem_reg_b3_b_b18_b (.CK(clk_i), .D(n_9347), .Q(u4_mem_b3_b_139), .SO(u4_mem_b3_b_139), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_138));
SDFFN u4_mem_reg_b3_b_b19_b (.CK(clk_i), .D(n_9345), .Q(u4_mem_b3_b_140), .SO(u4_mem_b3_b_140), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_139));
SDFFN u4_mem_reg_b3_b_b1_b (.CK(clk_i), .D(n_9344), .Q(u4_mem_b3_b_122), .SO(u4_mem_b3_b_122), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_140));
SDFFN u4_mem_reg_b3_b_b20_b (.CK(clk_i), .D(n_9343), .Q(u4_mem_b3_b_141), .SO(u4_mem_b3_b_141), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_122));
SDFFN u4_mem_reg_b3_b_b21_b (.CK(clk_i), .D(n_9342), .Q(u4_mem_b3_b_142), .SO(u4_mem_b3_b_142), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_141));
SDFFN u4_mem_reg_b3_b_b22_b (.CK(clk_i), .D(n_9340), .Q(u4_mem_b3_b_143), .SO(u4_mem_b3_b_143), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_142));
SDFFN u4_mem_reg_b3_b_b24_b (.CK(clk_i), .D(n_9338), .Q(u4_mem_b3_b_145), .SO(u4_mem_b3_b_145), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_143));
SDFFN u4_mem_reg_b3_b_b25_b (.CK(clk_i), .D(n_9337), .Q(u4_mem_b3_b_146), .SO(u4_mem_b3_b_146), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_145));
SDFFN u4_mem_reg_b3_b_b26_b (.CK(clk_i), .D(n_9335), .Q(u4_mem_b3_b_147), .SO(u4_mem_b3_b_147), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_146));
SDFFN u4_mem_reg_b3_b_b28_b (.CK(clk_i), .D(n_9332), .Q(u4_mem_b3_b_149), .SO(u4_mem_b3_b_149), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_147));
SDFFN u4_mem_reg_b3_b_b29_b (.CK(clk_i), .D(n_9331), .Q(u4_mem_b3_b_150), .SO(u4_mem_b3_b_150), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_149));
SDFFN u4_mem_reg_b3_b_b2_b (.CK(clk_i), .D(n_9330), .Q(u4_mem_b3_b_123), .SO(u4_mem_b3_b_123), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_150));
SDFFN u4_mem_reg_b3_b_b31_b (.CK(clk_i), .D(n_9328), .Q(u4_mem_b3_b_152), .SO(u4_mem_b3_b_152), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_123));
SDFFN u4_mem_reg_b3_b_b3_b (.CK(clk_i), .D(n_9327), .Q(u4_mem_b3_b_124), .SO(u4_mem_b3_b_124), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_152));
SDFFN u4_mem_reg_b3_b_b4_b (.CK(clk_i), .D(n_9325), .Q(u4_mem_b3_b_125), .SO(u4_mem_b3_b_125), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_124));
SDFFN u4_mem_reg_b3_b_b6_b (.CK(clk_i), .D(n_9322), .Q(u4_mem_b3_b_127), .SO(u4_mem_b3_b_127), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_125));
SDFFN u4_mem_reg_b3_b_b7_b (.CK(clk_i), .D(n_9321), .Q(u4_mem_b3_b_128), .SO(u4_mem_b3_b_128), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_127));
SDFFN u4_mem_reg_b3_b_b8_b (.CK(clk_i), .D(n_9320), .Q(u4_mem_b3_b_129), .SO(u4_mem_b3_b_129), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_128));
SDFFN u3_mem_reg_b2_b_b20_b (.CK(clk_i), .D(n_9195), .Q(u3_mem_b2_b_48), .SO(u3_mem_b2_b_48), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b3_b_129));
SDFFN u5_mem_reg_b1_b_b0_b (.CK(clk_i), .D(n_9317), .Q(u5_mem_b1_b), .SO(u5_mem_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b2_b_48));
SDFFN u5_mem_reg_b1_b_b10_b (.CK(clk_i), .D(n_9316), .Q(u5_mem_b1_b_69), .SO(u5_mem_b1_b_69), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b));
SDFFN u5_mem_reg_b1_b_b12_b (.CK(clk_i), .D(n_9314), .Q(u5_mem_b1_b_71), .SO(u5_mem_b1_b_71), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_69));
SDFFN u5_mem_reg_b1_b_b13_b (.CK(clk_i), .D(n_9313), .Q(u5_mem_b1_b_72), .SO(u5_mem_b1_b_72), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_71));
SDFFN u5_mem_reg_b1_b_b14_b (.CK(clk_i), .D(n_9312), .Q(u5_mem_b1_b_73), .SO(u5_mem_b1_b_73), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_72));
SDFFN u7_mem_reg_b1_b_b14_b (.CK(clk_i), .D(n_9060), .Q(u7_mem_b1_b_73), .SO(u7_mem_b1_b_73), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_73));
SDFFN u5_mem_reg_b1_b_b16_b (.CK(clk_i), .D(n_9308), .Q(u5_mem_b1_b_75), .SO(u5_mem_b1_b_75), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_73));
SDFFN u5_mem_reg_b1_b_b17_b (.CK(clk_i), .D(n_9306), .Q(u5_mem_b1_b_76), .SO(u5_mem_b1_b_76), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_75));
SDFFN u5_mem_reg_b1_b_b18_b (.CK(clk_i), .D(n_9304), .Q(u5_mem_b1_b_77), .SO(u5_mem_b1_b_77), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_76));
SDFFN u5_mem_reg_b1_b_b1_b (.CK(clk_i), .D(n_9301), .Q(u5_mem_b1_b_60), .SO(u5_mem_b1_b_60), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_77));
SDFFN u5_mem_reg_b1_b_b20_b (.CK(clk_i), .D(n_9300), .Q(u5_mem_b1_b_79), .SO(u5_mem_b1_b_79), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_60));
SDFFN u5_mem_reg_b1_b_b21_b (.CK(clk_i), .D(n_9299), .Q(u5_mem_b1_b_80), .SO(u5_mem_b1_b_80), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_79));
SDFFN u5_mem_reg_b1_b_b23_b (.CK(clk_i), .D(n_9297), .Q(u5_mem_b1_b_82), .SO(u5_mem_b1_b_82), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_80));
SDFFN u5_mem_reg_b1_b_b24_b (.CK(clk_i), .D(n_9296), .Q(u5_mem_b1_b_83), .SO(u5_mem_b1_b_83), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_82));
SDFFN u5_mem_reg_b1_b_b25_b (.CK(clk_i), .D(n_9294), .Q(u5_mem_b1_b_84), .SO(u5_mem_b1_b_84), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_83));
SDFFN u5_mem_reg_b1_b_b27_b (.CK(clk_i), .D(n_9292), .Q(u5_mem_b1_b_86), .SO(u5_mem_b1_b_86), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_84));
SDFFN u5_mem_reg_b1_b_b28_b (.CK(clk_i), .D(n_9291), .Q(u5_mem_b1_b_87), .SO(u5_mem_b1_b_87), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_86));
SDFFN u5_mem_reg_b1_b_b29_b (.CK(clk_i), .D(n_9289), .Q(u5_mem_b1_b_88), .SO(u5_mem_b1_b_88), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_87));
SDFFN u5_mem_reg_b1_b_b30_b (.CK(clk_i), .D(n_9285), .Q(u5_mem_b1_b_89), .SO(u5_mem_b1_b_89), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_88));
SDFFN u5_mem_reg_b1_b_b31_b (.CK(clk_i), .D(n_9283), .Q(u5_mem_b1_b_90), .SO(u5_mem_b1_b_90), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_89));
SDFFN u5_mem_reg_b1_b_b3_b (.CK(clk_i), .D(n_9282), .Q(u5_mem_b1_b_62), .SO(u5_mem_b1_b_62), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_90));
SDFFN u5_mem_reg_b1_b_b5_b (.CK(clk_i), .D(n_9280), .Q(u5_mem_b1_b_64), .SO(u5_mem_b1_b_64), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_62));
SDFFN u5_mem_reg_b1_b_b6_b (.CK(clk_i), .D(n_9278), .Q(u5_mem_b1_b_65), .SO(u5_mem_b1_b_65), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_64));
SDFFN u5_mem_reg_b1_b_b7_b (.CK(clk_i), .D(n_9277), .Q(u5_mem_b1_b_66), .SO(u5_mem_b1_b_66), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_65));
SDFFN u5_mem_reg_b1_b_b9_b (.CK(clk_i), .D(n_9275), .Q(u5_mem_b1_b_68), .SO(u5_mem_b1_b_68), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_66));
SDFFN u5_mem_reg_b2_b_b0_b (.CK(clk_i), .D(n_9274), .Q(u5_mem_b2_b), .SO(u5_mem_b2_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_68));
SDFFN u5_mem_reg_b2_b_b10_b (.CK(clk_i), .D(n_9273), .Q(u5_mem_b2_b_38), .SO(u5_mem_b2_b_38), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b));
SDFFN u5_mem_reg_b2_b_b12_b (.CK(clk_i), .D(n_9270), .Q(u5_mem_b2_b_40), .SO(u5_mem_b2_b_40), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_38));
SDFFN u5_mem_reg_b2_b_b13_b (.CK(clk_i), .D(n_9269), .Q(u5_mem_b2_b_41), .SO(u5_mem_b2_b_41), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_40));
SDFFN u5_mem_reg_b2_b_b14_b (.CK(clk_i), .D(n_9268), .Q(u5_mem_b2_b_42), .SO(u5_mem_b2_b_42), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_41));
SDFFN u5_mem_reg_b2_b_b16_b (.CK(clk_i), .D(n_9266), .Q(u5_mem_b2_b_44), .SO(u5_mem_b2_b_44), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_42));
SDFFN u5_mem_reg_b2_b_b17_b (.CK(clk_i), .D(n_9265), .Q(u5_mem_b2_b_45), .SO(u5_mem_b2_b_45), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_44));
SDFFN u5_mem_reg_b2_b_b18_b (.CK(clk_i), .D(n_9263), .Q(u5_mem_b2_b_46), .SO(u5_mem_b2_b_46), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_45));
SDFFN u5_mem_reg_b2_b_b1_b (.CK(clk_i), .D(n_9261), .Q(u5_mem_b2_b_29), .SO(u5_mem_b2_b_29), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_46));
SDFFN u5_mem_reg_b2_b_b20_b (.CK(clk_i), .D(n_9259), .Q(u5_mem_b2_b_48), .SO(u5_mem_b2_b_48), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_29));
SDFFN u5_mem_reg_b2_b_b21_b (.CK(clk_i), .D(n_9258), .Q(u5_mem_b2_b_49), .SO(u5_mem_b2_b_49), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_48));
SDFFN u5_mem_reg_b2_b_b23_b (.CK(clk_i), .D(n_9256), .Q(u5_mem_b2_b_51), .SO(u5_mem_b2_b_51), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_49));
SDFFN u5_mem_reg_b2_b_b24_b (.CK(clk_i), .D(n_9255), .Q(u5_mem_b2_b_52), .SO(u5_mem_b2_b_52), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_51));
SDFFN u5_mem_reg_b2_b_b25_b (.CK(clk_i), .D(n_9254), .Q(u5_mem_b2_b_53), .SO(u5_mem_b2_b_53), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_52));
SDFFN u5_mem_reg_b2_b_b27_b (.CK(clk_i), .D(n_9252), .Q(u5_mem_b2_b_55), .SO(u5_mem_b2_b_55), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_53));
SDFFN u5_mem_reg_b2_b_b28_b (.CK(clk_i), .D(n_9250), .Q(u5_mem_b2_b_56), .SO(u5_mem_b2_b_56), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_55));
SDFFN u5_mem_reg_b2_b_b29_b (.CK(clk_i), .D(n_9249), .Q(u5_mem_b2_b_57), .SO(u5_mem_b2_b_57), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_56));
SDFFN u5_mem_reg_b2_b_b30_b (.CK(clk_i), .D(n_9246), .Q(u5_mem_b2_b_58), .SO(u5_mem_b2_b_58), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_57));
SDFFN u5_mem_reg_b2_b_b31_b (.CK(clk_i), .D(n_9245), .Q(u5_mem_b2_b_59), .SO(u5_mem_b2_b_59), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_58));
SDFFN u5_mem_reg_b2_b_b3_b (.CK(clk_i), .D(n_9244), .Q(u5_mem_b2_b_31), .SO(u5_mem_b2_b_31), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_59));
SDFFN u5_mem_reg_b2_b_b4_b (.CK(clk_i), .D(n_9243), .Q(u5_mem_b2_b_32), .SO(u5_mem_b2_b_32), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_31));
SDFFN u5_mem_reg_b2_b_b5_b (.CK(clk_i), .D(n_9242), .Q(u5_mem_b2_b_33), .SO(u5_mem_b2_b_33), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_32));
SDFFN u5_mem_reg_b2_b_b6_b (.CK(clk_i), .D(n_9241), .Q(u5_mem_b2_b_34), .SO(u5_mem_b2_b_34), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_33));
SDFFN u5_mem_reg_b2_b_b7_b (.CK(clk_i), .D(n_9240), .Q(u5_mem_b2_b_35), .SO(u5_mem_b2_b_35), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_34));
SDFFN u5_mem_reg_b2_b_b9_b (.CK(clk_i), .D(n_9238), .Q(u5_mem_b2_b_37), .SO(u5_mem_b2_b_37), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_35));
SDFFN u5_mem_reg_b3_b_b0_b (.CK(clk_i), .D(n_9237), .Q(u5_mem_b3_b), .SO(u5_mem_b3_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_37));
SDFFN u5_mem_reg_b3_b_b10_b (.CK(clk_i), .D(n_9236), .Q(u5_mem_b3_b_131), .SO(u5_mem_b3_b_131), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b));
SDFFN u5_mem_reg_b3_b_b12_b (.CK(clk_i), .D(n_9233), .Q(u5_mem_b3_b_133), .SO(u5_mem_b3_b_133), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_131));
SDFFN u5_mem_reg_b3_b_b13_b (.CK(clk_i), .D(n_9232), .Q(u5_mem_b3_b_134), .SO(u5_mem_b3_b_134), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_133));
SDFFN u5_mem_reg_b3_b_b14_b (.CK(clk_i), .D(n_9231), .Q(u5_mem_b3_b_135), .SO(u5_mem_b3_b_135), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_134));
SDFFN u5_mem_reg_b3_b_b16_b (.CK(clk_i), .D(n_9228), .Q(u5_mem_b3_b_137), .SO(u5_mem_b3_b_137), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_135));
SDFFN u5_mem_reg_b3_b_b17_b (.CK(clk_i), .D(n_9227), .Q(u5_mem_b3_b_138), .SO(u5_mem_b3_b_138), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_137));
SDFFN u5_mem_reg_b3_b_b18_b (.CK(clk_i), .D(n_9226), .Q(u5_mem_b3_b_139), .SO(u5_mem_b3_b_139), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_138));
SDFFN u5_mem_reg_b3_b_b1_b (.CK(clk_i), .D(n_9223), .Q(u5_mem_b3_b_122), .SO(u5_mem_b3_b_122), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_139));
SDFFN u5_mem_reg_b3_b_b20_b (.CK(clk_i), .D(n_9222), .Q(u5_mem_b3_b_141), .SO(u5_mem_b3_b_141), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_122));
SDFFN u5_mem_reg_b3_b_b21_b (.CK(clk_i), .D(n_9221), .Q(u5_mem_b3_b_142), .SO(u5_mem_b3_b_142), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_141));
SDFFN u6_mem_reg_b0_b_b17_b (.CK(clk_i), .D(n_8775), .Q(u6_mem_b0_b_107), .SO(u6_mem_b0_b_107), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_142));
SDFFN u5_mem_reg_b3_b_b23_b (.CK(clk_i), .D(n_9218), .Q(u5_mem_b3_b_144), .SO(u5_mem_b3_b_144), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_107));
SDFFN u5_mem_reg_b3_b_b24_b (.CK(clk_i), .D(n_9217), .Q(u5_mem_b3_b_145), .SO(u5_mem_b3_b_145), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_144));
SDFFN u5_mem_reg_b3_b_b25_b (.CK(clk_i), .D(n_9216), .Q(u5_mem_b3_b_146), .SO(u5_mem_b3_b_146), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_145));
SDFFN u5_mem_reg_b3_b_b27_b (.CK(clk_i), .D(n_9213), .Q(u5_mem_b3_b_148), .SO(u5_mem_b3_b_148), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_146));
SDFFN u5_mem_reg_b3_b_b28_b (.CK(clk_i), .D(n_9211), .Q(u5_mem_b3_b_149), .SO(u5_mem_b3_b_149), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_148));
SDFFN u5_mem_reg_b3_b_b29_b (.CK(clk_i), .D(n_9210), .Q(u5_mem_b3_b_150), .SO(u5_mem_b3_b_150), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_149));
SDFFN u5_mem_reg_b3_b_b30_b (.CK(clk_i), .D(n_9208), .Q(u5_mem_b3_b_151), .SO(u5_mem_b3_b_151), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_150));
SDFFN u5_mem_reg_b3_b_b31_b (.CK(clk_i), .D(n_9207), .Q(u5_mem_b3_b_152), .SO(u5_mem_b3_b_152), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_151));
SDFFN u5_mem_reg_b3_b_b3_b (.CK(clk_i), .D(n_9206), .Q(u5_mem_b3_b_124), .SO(u5_mem_b3_b_124), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_152));
SDFFN u5_mem_reg_b3_b_b5_b (.CK(clk_i), .D(n_9203), .Q(u5_mem_b3_b_126), .SO(u5_mem_b3_b_126), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_124));
SDFFN u5_mem_reg_b3_b_b6_b (.CK(clk_i), .D(n_9201), .Q(u5_mem_b3_b_127), .SO(u5_mem_b3_b_127), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_126));
SDFFN u5_mem_reg_b3_b_b7_b (.CK(clk_i), .D(n_9200), .Q(u5_mem_b3_b_128), .SO(u5_mem_b3_b_128), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_127));
SDFFN u5_mem_reg_b3_b_b9_b (.CK(clk_i), .D(n_9198), .Q(u5_mem_b3_b_130), .SO(u5_mem_b3_b_130), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_128));
SDFFN u6_mem_reg_b1_b_b0_b (.CK(clk_i), .D(n_9192), .Q(u6_mem_b1_b), .SO(u6_mem_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_130));
SDFFN u6_mem_reg_b1_b_b10_b (.CK(clk_i), .D(n_9191), .Q(u6_mem_b1_b_69), .SO(u6_mem_b1_b_69), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b));
SDFFN u6_mem_reg_b1_b_b12_b (.CK(clk_i), .D(n_9189), .Q(u6_mem_b1_b_71), .SO(u6_mem_b1_b_71), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_69));
SDFFN u6_mem_reg_b1_b_b13_b (.CK(clk_i), .D(n_9188), .Q(u6_mem_b1_b_72), .SO(u6_mem_b1_b_72), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_71));
SDFFN u6_mem_reg_b1_b_b14_b (.CK(clk_i), .D(n_9187), .Q(u6_mem_b1_b_73), .SO(u6_mem_b1_b_73), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_72));
SDFFN u6_mem_reg_b1_b_b16_b (.CK(clk_i), .D(n_9183), .Q(u6_mem_b1_b_75), .SO(u6_mem_b1_b_75), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_73));
SDFFN u6_mem_reg_b1_b_b17_b (.CK(clk_i), .D(n_9181), .Q(u6_mem_b1_b_76), .SO(u6_mem_b1_b_76), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_75));
SDFFN u6_mem_reg_b1_b_b18_b (.CK(clk_i), .D(n_9179), .Q(u6_mem_b1_b_77), .SO(u6_mem_b1_b_77), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_76));
SDFFN u6_mem_reg_b1_b_b19_b (.CK(clk_i), .D(n_9177), .Q(u6_mem_b1_b_78), .SO(u6_mem_b1_b_78), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_77));
SDFFN u6_mem_reg_b1_b_b1_b (.CK(clk_i), .D(n_9176), .Q(u6_mem_b1_b_60), .SO(u6_mem_b1_b_60), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_78));
SDFFN u6_mem_reg_b1_b_b20_b (.CK(clk_i), .D(n_9175), .Q(u6_mem_b1_b_79), .SO(u6_mem_b1_b_79), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_60));
SDFFN u6_mem_reg_b1_b_b21_b (.CK(clk_i), .D(n_9174), .Q(u6_mem_b1_b_80), .SO(u6_mem_b1_b_80), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_79));
SDFFN u6_mem_reg_b1_b_b23_b (.CK(clk_i), .D(n_9172), .Q(u6_mem_b1_b_82), .SO(u6_mem_b1_b_82), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_80));
SDFFN u6_mem_reg_b1_b_b24_b (.CK(clk_i), .D(n_9171), .Q(u6_mem_b1_b_83), .SO(u6_mem_b1_b_83), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_82));
SDFFN u6_mem_reg_b1_b_b25_b (.CK(clk_i), .D(n_9169), .Q(u6_mem_b1_b_84), .SO(u6_mem_b1_b_84), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_83));
SDFFN u6_mem_reg_b1_b_b27_b (.CK(clk_i), .D(n_9167), .Q(u6_mem_b1_b_86), .SO(u6_mem_b1_b_86), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_84));
SDFFN u6_mem_reg_b1_b_b28_b (.CK(clk_i), .D(n_9166), .Q(u6_mem_b1_b_87), .SO(u6_mem_b1_b_87), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_86));
SDFFN u6_mem_reg_b1_b_b29_b (.CK(clk_i), .D(n_9164), .Q(u6_mem_b1_b_88), .SO(u6_mem_b1_b_88), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_87));
SDFFN u6_mem_reg_b1_b_b30_b (.CK(clk_i), .D(n_9160), .Q(u6_mem_b1_b_89), .SO(u6_mem_b1_b_89), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_88));
SDFFN u6_mem_reg_b1_b_b31_b (.CK(clk_i), .D(n_9158), .Q(u6_mem_b1_b_90), .SO(u6_mem_b1_b_90), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_89));
SDFFN u6_mem_reg_b1_b_b3_b (.CK(clk_i), .D(n_9157), .Q(u6_mem_b1_b_62), .SO(u6_mem_b1_b_62), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_90));
SDFFN u6_mem_reg_b1_b_b5_b (.CK(clk_i), .D(n_9155), .Q(u6_mem_b1_b_64), .SO(u6_mem_b1_b_64), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_62));
SDFFN u6_mem_reg_b1_b_b6_b (.CK(clk_i), .D(n_9153), .Q(u6_mem_b1_b_65), .SO(u6_mem_b1_b_65), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_64));
SDFFN u6_mem_reg_b1_b_b7_b (.CK(clk_i), .D(n_9152), .Q(u6_mem_b1_b_66), .SO(u6_mem_b1_b_66), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_65));
SDFFN u6_mem_reg_b1_b_b9_b (.CK(clk_i), .D(n_9150), .Q(u6_mem_b1_b_68), .SO(u6_mem_b1_b_68), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_66));
SDFFN u6_mem_reg_b2_b_b0_b (.CK(clk_i), .D(n_9149), .Q(u6_mem_b2_b), .SO(u6_mem_b2_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_68));
SDFFN u6_mem_reg_b2_b_b10_b (.CK(clk_i), .D(n_9148), .Q(u6_mem_b2_b_38), .SO(u6_mem_b2_b_38), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b));
SDFFN u6_mem_reg_b2_b_b12_b (.CK(clk_i), .D(n_9145), .Q(u6_mem_b2_b_40), .SO(u6_mem_b2_b_40), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_38));
SDFFN u6_mem_reg_b2_b_b13_b (.CK(clk_i), .D(n_9144), .Q(u6_mem_b2_b_41), .SO(u6_mem_b2_b_41), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_40));
SDFFN u6_mem_reg_b2_b_b14_b (.CK(clk_i), .D(n_9143), .Q(u6_mem_b2_b_42), .SO(u6_mem_b2_b_42), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_41));
SDFFN u6_mem_reg_b2_b_b16_b (.CK(clk_i), .D(n_9141), .Q(u6_mem_b2_b_44), .SO(u6_mem_b2_b_44), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_42));
SDFFN u6_mem_reg_b2_b_b17_b (.CK(clk_i), .D(n_9140), .Q(u6_mem_b2_b_45), .SO(u6_mem_b2_b_45), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_44));
SDFFN u6_mem_reg_b2_b_b18_b (.CK(clk_i), .D(n_9138), .Q(u6_mem_b2_b_46), .SO(u6_mem_b2_b_46), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_45));
SDFFN u6_mem_reg_b2_b_b1_b (.CK(clk_i), .D(n_9136), .Q(u6_mem_b2_b_29), .SO(u6_mem_b2_b_29), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_46));
SDFFN u6_mem_reg_b2_b_b20_b (.CK(clk_i), .D(n_9134), .Q(u6_mem_b2_b_48), .SO(u6_mem_b2_b_48), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_29));
SDFFN u6_mem_reg_b2_b_b21_b (.CK(clk_i), .D(n_9133), .Q(u6_mem_b2_b_49), .SO(u6_mem_b2_b_49), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_48));
SDFFN u6_mem_reg_b2_b_b23_b (.CK(clk_i), .D(n_9131), .Q(u6_mem_b2_b_51), .SO(u6_mem_b2_b_51), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_49));
SDFFN u6_mem_reg_b2_b_b24_b (.CK(clk_i), .D(n_9130), .Q(u6_mem_b2_b_52), .SO(u6_mem_b2_b_52), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_51));
SDFFN u6_mem_reg_b2_b_b25_b (.CK(clk_i), .D(n_9129), .Q(u6_mem_b2_b_53), .SO(u6_mem_b2_b_53), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_52));
SDFFN u6_mem_reg_b2_b_b27_b (.CK(clk_i), .D(n_9127), .Q(u6_mem_b2_b_55), .SO(u6_mem_b2_b_55), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_53));
SDFFN u6_mem_reg_b2_b_b28_b (.CK(clk_i), .D(n_9125), .Q(u6_mem_b2_b_56), .SO(u6_mem_b2_b_56), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_55));
SDFFN u6_mem_reg_b2_b_b29_b (.CK(clk_i), .D(n_9124), .Q(u6_mem_b2_b_57), .SO(u6_mem_b2_b_57), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_56));
SDFFN u6_mem_reg_b2_b_b30_b (.CK(clk_i), .D(n_9121), .Q(u6_mem_b2_b_58), .SO(u6_mem_b2_b_58), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_57));
SDFFN u6_mem_reg_b2_b_b31_b (.CK(clk_i), .D(n_9120), .Q(u6_mem_b2_b_59), .SO(u6_mem_b2_b_59), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_58));
SDFFN u6_mem_reg_b2_b_b3_b (.CK(clk_i), .D(n_9119), .Q(u6_mem_b2_b_31), .SO(u6_mem_b2_b_31), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_59));
SDFFN u6_mem_reg_b2_b_b5_b (.CK(clk_i), .D(n_9117), .Q(u6_mem_b2_b_33), .SO(u6_mem_b2_b_33), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_31));
SDFFN u6_mem_reg_b2_b_b6_b (.CK(clk_i), .D(n_9116), .Q(u6_mem_b2_b_34), .SO(u6_mem_b2_b_34), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_33));
SDFFN u6_mem_reg_b2_b_b7_b (.CK(clk_i), .D(n_9115), .Q(u6_mem_b2_b_35), .SO(u6_mem_b2_b_35), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_34));
SDFFN u6_mem_reg_b2_b_b9_b (.CK(clk_i), .D(n_9113), .Q(u6_mem_b2_b_37), .SO(u6_mem_b2_b_37), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_35));
SDFFN u6_mem_reg_b3_b_b0_b (.CK(clk_i), .D(n_9112), .Q(u6_mem_b3_b), .SO(u6_mem_b3_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_37));
SDFFN u6_mem_reg_b3_b_b10_b (.CK(clk_i), .D(n_9111), .Q(u6_mem_b3_b_131), .SO(u6_mem_b3_b_131), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b));
SDFFN u6_mem_reg_b3_b_b12_b (.CK(clk_i), .D(n_9108), .Q(u6_mem_b3_b_133), .SO(u6_mem_b3_b_133), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_131));
SDFFN u6_mem_reg_b3_b_b13_b (.CK(clk_i), .D(n_9107), .Q(u6_mem_b3_b_134), .SO(u6_mem_b3_b_134), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_133));
SDFFN u6_mem_reg_b3_b_b14_b (.CK(clk_i), .D(n_9106), .Q(u6_mem_b3_b_135), .SO(u6_mem_b3_b_135), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_134));
SDFFN u6_mem_reg_b3_b_b16_b (.CK(clk_i), .D(n_9103), .Q(u6_mem_b3_b_137), .SO(u6_mem_b3_b_137), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_135));
SDFFN u6_mem_reg_b3_b_b17_b (.CK(clk_i), .D(n_9102), .Q(u6_mem_b3_b_138), .SO(u6_mem_b3_b_138), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_137));
SDFFN u6_mem_reg_b3_b_b18_b (.CK(clk_i), .D(n_9101), .Q(u6_mem_b3_b_139), .SO(u6_mem_b3_b_139), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_138));
SDFFN u6_mem_reg_b3_b_b1_b (.CK(clk_i), .D(n_9098), .Q(u6_mem_b3_b_122), .SO(u6_mem_b3_b_122), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_139));
SDFFN u6_mem_reg_b3_b_b20_b (.CK(clk_i), .D(n_9097), .Q(u6_mem_b3_b_141), .SO(u6_mem_b3_b_141), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_122));
SDFFN u6_mem_reg_b3_b_b21_b (.CK(clk_i), .D(n_9096), .Q(u6_mem_b3_b_142), .SO(u6_mem_b3_b_142), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_141));
SDFFN u6_mem_reg_b3_b_b23_b (.CK(clk_i), .D(n_9093), .Q(u6_mem_b3_b_144), .SO(u6_mem_b3_b_144), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_142));
SDFFN u6_mem_reg_b3_b_b24_b (.CK(clk_i), .D(n_9092), .Q(u6_mem_b3_b_145), .SO(u6_mem_b3_b_145), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_144));
SDFFN u6_mem_reg_b3_b_b25_b (.CK(clk_i), .D(n_9091), .Q(u6_mem_b3_b_146), .SO(u6_mem_b3_b_146), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_145));
SDFFN u6_mem_reg_b3_b_b27_b (.CK(clk_i), .D(n_9088), .Q(u6_mem_b3_b_148), .SO(u6_mem_b3_b_148), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_146));
SDFFN u6_mem_reg_b3_b_b28_b (.CK(clk_i), .D(n_9086), .Q(u6_mem_b3_b_149), .SO(u6_mem_b3_b_149), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_148));
SDFFN u6_mem_reg_b3_b_b29_b (.CK(clk_i), .D(n_9085), .Q(u6_mem_b3_b_150), .SO(u6_mem_b3_b_150), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_149));
SDFFN u6_mem_reg_b3_b_b30_b (.CK(clk_i), .D(n_9083), .Q(u6_mem_b3_b_151), .SO(u6_mem_b3_b_151), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_150));
SDFFN u6_mem_reg_b3_b_b31_b (.CK(clk_i), .D(n_9082), .Q(u6_mem_b3_b_152), .SO(u6_mem_b3_b_152), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_151));
SDFFN u6_mem_reg_b3_b_b3_b (.CK(clk_i), .D(n_9081), .Q(u6_mem_b3_b_124), .SO(u6_mem_b3_b_124), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_152));
SDFFN u6_mem_reg_b3_b_b5_b (.CK(clk_i), .D(n_9078), .Q(u6_mem_b3_b_126), .SO(u6_mem_b3_b_126), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_124));
SDFFN u6_mem_reg_b3_b_b6_b (.CK(clk_i), .D(n_9076), .Q(u6_mem_b3_b_127), .SO(u6_mem_b3_b_127), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_126));
SDFFN u6_mem_reg_b3_b_b7_b (.CK(clk_i), .D(n_9075), .Q(u6_mem_b3_b_128), .SO(u6_mem_b3_b_128), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_127));
SDFFN u6_mem_reg_b3_b_b9_b (.CK(clk_i), .D(n_9073), .Q(u6_mem_b3_b_130), .SO(u6_mem_b3_b_130), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_128));
SDFFN u3_mem_reg_b3_b_b8_b (.CK(clk_i), .D(n_8353), .Q(u3_mem_b3_b_129), .SO(u3_mem_b3_b_129), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_130));
SDFFN u7_mem_reg_b1_b_b0_b (.CK(clk_i), .D(n_9066), .Q(u7_mem_b1_b), .SO(u7_mem_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b3_b_129));
SDFFN u7_mem_reg_b1_b_b11_b (.CK(clk_i), .D(n_9064), .Q(u7_mem_b1_b_70), .SO(u7_mem_b1_b_70), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b));
SDFFN u7_mem_reg_b1_b_b12_b (.CK(clk_i), .D(n_9062), .Q(u7_mem_b1_b_71), .SO(u7_mem_b1_b_71), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_70));
SDFFN u7_mem_reg_b1_b_b13_b (.CK(clk_i), .D(n_9061), .Q(u7_mem_b1_b_72), .SO(u7_mem_b1_b_72), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_71));
SDFFN u7_mem_reg_b1_b_b15_b (.CK(clk_i), .D(n_9058), .Q(u7_mem_b1_b_74), .SO(u7_mem_b1_b_74), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_72));
SDFFN u7_mem_reg_b1_b_b16_b (.CK(clk_i), .D(n_9056), .Q(u7_mem_b1_b_75), .SO(u7_mem_b1_b_75), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_74));
SDFFN u7_mem_reg_b1_b_b17_b (.CK(clk_i), .D(n_9054), .Q(u7_mem_b1_b_76), .SO(u7_mem_b1_b_76), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_75));
SDFFN u7_mem_reg_b1_b_b18_b (.CK(clk_i), .D(n_9052), .Q(u7_mem_b1_b_77), .SO(u7_mem_b1_b_77), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_76));
SDFFN u7_mem_reg_b1_b_b19_b (.CK(clk_i), .D(n_9050), .Q(u7_mem_b1_b_78), .SO(u7_mem_b1_b_78), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_77));
SDFFN u7_mem_reg_b1_b_b1_b (.CK(clk_i), .D(n_9049), .Q(u7_mem_b1_b_60), .SO(u7_mem_b1_b_60), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_78));
SDFFN u7_mem_reg_b1_b_b20_b (.CK(clk_i), .D(n_9048), .Q(u7_mem_b1_b_79), .SO(u7_mem_b1_b_79), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_60));
SDFFN u7_mem_reg_b1_b_b22_b (.CK(clk_i), .D(n_9046), .Q(u7_mem_b1_b_81), .SO(u7_mem_b1_b_81), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_79));
SDFFN u7_mem_reg_b1_b_b23_b (.CK(clk_i), .D(n_9045), .Q(u7_mem_b1_b_82), .SO(u7_mem_b1_b_82), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_81));
SDFFN u7_mem_reg_b1_b_b24_b (.CK(clk_i), .D(n_9044), .Q(u7_mem_b1_b_83), .SO(u7_mem_b1_b_83), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_82));
SDFFN u7_mem_reg_b1_b_b26_b (.CK(clk_i), .D(n_9041), .Q(u7_mem_b1_b_85), .SO(u7_mem_b1_b_85), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_83));
SDFFN u7_mem_reg_b1_b_b27_b (.CK(clk_i), .D(n_9040), .Q(u7_mem_b1_b_86), .SO(u7_mem_b1_b_86), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_85));
SDFFN u7_mem_reg_b1_b_b28_b (.CK(clk_i), .D(n_9039), .Q(u7_mem_b1_b_87), .SO(u7_mem_b1_b_87), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_86));
SDFFN u7_mem_reg_b1_b_b2_b (.CK(clk_i), .D(n_9035), .Q(u7_mem_b1_b_61), .SO(u7_mem_b1_b_61), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_87));
SDFFN u7_mem_reg_b1_b_b30_b (.CK(clk_i), .D(n_9033), .Q(u7_mem_b1_b_89), .SO(u7_mem_b1_b_89), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_61));
SDFFN u7_mem_reg_b1_b_b31_b (.CK(clk_i), .D(n_9031), .Q(u7_mem_b1_b_90), .SO(u7_mem_b1_b_90), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_89));
SDFFN u7_mem_reg_b1_b_b4_b (.CK(clk_i), .D(n_9029), .Q(u7_mem_b1_b_63), .SO(u7_mem_b1_b_63), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_90));
SDFFN u7_mem_reg_b1_b_b5_b (.CK(clk_i), .D(n_9028), .Q(u7_mem_b1_b_64), .SO(u7_mem_b1_b_64), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_63));
SDFFN u7_mem_reg_b1_b_b6_b (.CK(clk_i), .D(n_9026), .Q(u7_mem_b1_b_65), .SO(u7_mem_b1_b_65), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_64));
SDFFN u7_mem_reg_b1_b_b8_b (.CK(clk_i), .D(n_9024), .Q(u7_mem_b1_b_67), .SO(u7_mem_b1_b_67), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_65));
SDFFN u7_mem_reg_b1_b_b9_b (.CK(clk_i), .D(n_9021), .Q(u7_mem_b1_b_68), .SO(u7_mem_b1_b_68), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_67));
SDFFN u7_mem_reg_b2_b_b0_b (.CK(clk_i), .D(n_9020), .Q(u7_mem_b2_b), .SO(u7_mem_b2_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_68));
SDFFN u7_mem_reg_b2_b_b11_b (.CK(clk_i), .D(n_9018), .Q(u7_mem_b2_b_39), .SO(u7_mem_b2_b_39), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b));
SDFFN u7_mem_reg_b2_b_b12_b (.CK(clk_i), .D(n_9016), .Q(u7_mem_b2_b_40), .SO(u7_mem_b2_b_40), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_39));
SDFFN u7_mem_reg_b2_b_b13_b (.CK(clk_i), .D(n_9015), .Q(u7_mem_b2_b_41), .SO(u7_mem_b2_b_41), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_40));
SDFFN u7_mem_reg_b2_b_b15_b (.CK(clk_i), .D(n_9013), .Q(u7_mem_b2_b_43), .SO(u7_mem_b2_b_43), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_41));
SDFFN u7_mem_reg_b2_b_b16_b (.CK(clk_i), .D(n_9012), .Q(u7_mem_b2_b_44), .SO(u7_mem_b2_b_44), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_43));
SDFFN u7_mem_reg_b2_b_b17_b (.CK(clk_i), .D(n_9011), .Q(u7_mem_b2_b_45), .SO(u7_mem_b2_b_45), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_44));
SDFFN u7_mem_reg_b2_b_b19_b (.CK(clk_i), .D(n_9008), .Q(u7_mem_b2_b_47), .SO(u7_mem_b2_b_47), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_45));
SDFFN u7_mem_reg_b2_b_b1_b (.CK(clk_i), .D(n_9007), .Q(u7_mem_b2_b_29), .SO(u7_mem_b2_b_29), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_47));
SDFFN u7_mem_reg_b2_b_b20_b (.CK(clk_i), .D(n_9005), .Q(u7_mem_b2_b_48), .SO(u7_mem_b2_b_48), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_29));
SDFFN u7_mem_reg_b2_b_b22_b (.CK(clk_i), .D(n_9003), .Q(u7_mem_b2_b_50), .SO(u7_mem_b2_b_50), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_48));
SDFFN u7_mem_reg_b2_b_b23_b (.CK(clk_i), .D(n_9002), .Q(u7_mem_b2_b_51), .SO(u7_mem_b2_b_51), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_50));
SDFFN u7_mem_reg_b2_b_b24_b (.CK(clk_i), .D(n_9001), .Q(u7_mem_b2_b_52), .SO(u7_mem_b2_b_52), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_51));
SDFFN u7_mem_reg_b2_b_b26_b (.CK(clk_i), .D(n_8999), .Q(u7_mem_b2_b_54), .SO(u7_mem_b2_b_54), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_52));
SDFFN u7_mem_reg_b2_b_b27_b (.CK(clk_i), .D(n_8998), .Q(u7_mem_b2_b_55), .SO(u7_mem_b2_b_55), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_54));
SDFFN u7_mem_reg_b2_b_b28_b (.CK(clk_i), .D(n_8996), .Q(u7_mem_b2_b_56), .SO(u7_mem_b2_b_56), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_55));
SDFFN u7_mem_reg_b2_b_b2_b (.CK(clk_i), .D(n_8993), .Q(u7_mem_b2_b_30), .SO(u7_mem_b2_b_30), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_56));
SDFFN u7_mem_reg_b2_b_b30_b (.CK(clk_i), .D(n_8992), .Q(u7_mem_b2_b_58), .SO(u7_mem_b2_b_58), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_30));
SDFFN u7_mem_reg_b2_b_b31_b (.CK(clk_i), .D(n_8991), .Q(u7_mem_b2_b_59), .SO(u7_mem_b2_b_59), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_58));
SDFFN u7_mem_reg_b2_b_b4_b (.CK(clk_i), .D(n_8989), .Q(u7_mem_b2_b_32), .SO(u7_mem_b2_b_32), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_59));
SDFFN u7_mem_reg_b2_b_b5_b (.CK(clk_i), .D(n_8988), .Q(u7_mem_b2_b_33), .SO(u7_mem_b2_b_33), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_32));
SDFFN u7_mem_reg_b2_b_b6_b (.CK(clk_i), .D(n_8987), .Q(u7_mem_b2_b_34), .SO(u7_mem_b2_b_34), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_33));
SDFFN u7_mem_reg_b2_b_b8_b (.CK(clk_i), .D(n_8985), .Q(u7_mem_b2_b_36), .SO(u7_mem_b2_b_36), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_34));
SDFFN u7_mem_reg_b2_b_b9_b (.CK(clk_i), .D(n_8984), .Q(u7_mem_b2_b_37), .SO(u7_mem_b2_b_37), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_36));
SDFFN u7_mem_reg_b3_b_b0_b (.CK(clk_i), .D(n_8983), .Q(u7_mem_b3_b), .SO(u7_mem_b3_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b2_b_37));
SDFFN u7_mem_reg_b3_b_b11_b (.CK(clk_i), .D(n_8980), .Q(u7_mem_b3_b_132), .SO(u7_mem_b3_b_132), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b));
SDFFN u7_mem_reg_b3_b_b12_b (.CK(clk_i), .D(n_8979), .Q(u7_mem_b3_b_133), .SO(u7_mem_b3_b_133), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_132));
SDFFN u7_mem_reg_b3_b_b13_b (.CK(clk_i), .D(n_8978), .Q(u7_mem_b3_b_134), .SO(u7_mem_b3_b_134), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_133));
SDFFN u7_mem_reg_b3_b_b15_b (.CK(clk_i), .D(n_8975), .Q(u7_mem_b3_b_136), .SO(u7_mem_b3_b_136), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_134));
SDFFN u7_mem_reg_b3_b_b16_b (.CK(clk_i), .D(n_8974), .Q(u7_mem_b3_b_137), .SO(u7_mem_b3_b_137), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_136));
SDFFN u7_mem_reg_b3_b_b17_b (.CK(clk_i), .D(n_8973), .Q(u7_mem_b3_b_138), .SO(u7_mem_b3_b_138), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_137));
SDFFN u7_mem_reg_b3_b_b19_b (.CK(clk_i), .D(n_8970), .Q(u7_mem_b3_b_140), .SO(u7_mem_b3_b_140), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_138));
SDFFN u7_mem_reg_b3_b_b1_b (.CK(clk_i), .D(n_8969), .Q(u7_mem_b3_b_122), .SO(u7_mem_b3_b_122), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_140));
SDFFN u7_mem_reg_b3_b_b20_b (.CK(clk_i), .D(n_8968), .Q(u7_mem_b3_b_141), .SO(u7_mem_b3_b_141), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_122));
SDFFN u6_mem_reg_b0_b_b20_b (.CK(clk_i), .D(n_8770), .Q(u6_mem_b0_b_110), .SO(u6_mem_b0_b_110), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_141));
SDFFN u7_mem_reg_b3_b_b22_b (.CK(clk_i), .D(n_8965), .Q(u7_mem_b3_b_143), .SO(u7_mem_b3_b_143), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_110));
SDFFN u7_mem_reg_b3_b_b23_b (.CK(clk_i), .D(n_8964), .Q(u7_mem_b3_b_144), .SO(u7_mem_b3_b_144), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_143));
SDFFN u7_mem_reg_b3_b_b24_b (.CK(clk_i), .D(n_8963), .Q(u7_mem_b3_b_145), .SO(u7_mem_b3_b_145), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_144));
SDFFN u7_mem_reg_b3_b_b26_b (.CK(clk_i), .D(n_8960), .Q(u7_mem_b3_b_147), .SO(u7_mem_b3_b_147), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_145));
SDFFN u7_mem_reg_b3_b_b27_b (.CK(clk_i), .D(n_8959), .Q(u7_mem_b3_b_148), .SO(u7_mem_b3_b_148), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_147));
SDFFN u7_mem_reg_b3_b_b28_b (.CK(clk_i), .D(n_8957), .Q(u7_mem_b3_b_149), .SO(u7_mem_b3_b_149), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_148));
SDFFN u7_mem_reg_b3_b_b2_b (.CK(clk_i), .D(n_8955), .Q(u7_mem_b3_b_123), .SO(u7_mem_b3_b_123), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_149));
SDFFN u7_mem_reg_b3_b_b30_b (.CK(clk_i), .D(n_8954), .Q(u7_mem_b3_b_151), .SO(u7_mem_b3_b_151), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_123));
SDFFN u7_mem_reg_b3_b_b31_b (.CK(clk_i), .D(n_8953), .Q(u7_mem_b3_b_152), .SO(u7_mem_b3_b_152), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_151));
SDFFN u7_mem_reg_b3_b_b4_b (.CK(clk_i), .D(n_8950), .Q(u7_mem_b3_b_125), .SO(u7_mem_b3_b_125), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_152));
SDFFN u7_mem_reg_b3_b_b5_b (.CK(clk_i), .D(n_8949), .Q(u7_mem_b3_b_126), .SO(u7_mem_b3_b_126), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_125));
SDFFN u7_mem_reg_b3_b_b6_b (.CK(clk_i), .D(n_8947), .Q(u7_mem_b3_b_127), .SO(u7_mem_b3_b_127), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_126));
SDFFN u7_mem_reg_b3_b_b8_b (.CK(clk_i), .D(n_8945), .Q(u7_mem_b3_b_129), .SO(u7_mem_b3_b_129), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_127));
SDFFN u7_mem_reg_b3_b_b9_b (.CK(clk_i), .D(n_8944), .Q(u7_mem_b3_b_130), .SO(u7_mem_b3_b_130), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_129));
SDFFN u8_mem_reg_b1_b_b0_b (.CK(clk_i), .D(n_8941), .Q(u8_mem_b1_b), .SO(u8_mem_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b3_b_130));
SDFFN u8_mem_reg_b1_b_b11_b (.CK(clk_i), .D(n_8939), .Q(u8_mem_b1_b_70), .SO(u8_mem_b1_b_70), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b));
SDFFN u8_mem_reg_b1_b_b12_b (.CK(clk_i), .D(n_8938), .Q(u8_mem_b1_b_71), .SO(u8_mem_b1_b_71), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_70));
SDFFN u8_mem_reg_b1_b_b13_b (.CK(clk_i), .D(n_8936), .Q(u8_mem_b1_b_72), .SO(u8_mem_b1_b_72), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_71));
SDFFN u8_mem_reg_b1_b_b15_b (.CK(clk_i), .D(n_8934), .Q(u8_mem_b1_b_74), .SO(u8_mem_b1_b_74), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_72));
SDFFN u8_mem_reg_b1_b_b16_b (.CK(clk_i), .D(n_8932), .Q(u8_mem_b1_b_75), .SO(u8_mem_b1_b_75), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_74));
SDFFN u8_mem_reg_b1_b_b17_b (.CK(clk_i), .D(n_8931), .Q(u8_mem_b1_b_76), .SO(u8_mem_b1_b_76), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_75));
SDFFN u8_mem_reg_b1_b_b19_b (.CK(clk_i), .D(n_8928), .Q(u8_mem_b1_b_78), .SO(u8_mem_b1_b_78), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_76));
SDFFN u8_mem_reg_b1_b_b1_b (.CK(clk_i), .D(n_8926), .Q(u8_mem_b1_b_60), .SO(u8_mem_b1_b_60), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_78));
SDFFN u8_mem_reg_b1_b_b20_b (.CK(clk_i), .D(n_8925), .Q(u8_mem_b1_b_79), .SO(u8_mem_b1_b_79), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_60));
SDFFN u8_mem_reg_b1_b_b22_b (.CK(clk_i), .D(n_8922), .Q(u8_mem_b1_b_81), .SO(u8_mem_b1_b_81), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_79));
SDFFN u8_mem_reg_b1_b_b23_b (.CK(clk_i), .D(n_8921), .Q(u8_mem_b1_b_82), .SO(u8_mem_b1_b_82), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_81));
SDFFN u8_mem_reg_b1_b_b24_b (.CK(clk_i), .D(n_8920), .Q(u8_mem_b1_b_83), .SO(u8_mem_b1_b_83), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_82));
SDFFN u8_mem_reg_b1_b_b26_b (.CK(clk_i), .D(n_8916), .Q(u8_mem_b1_b_85), .SO(u8_mem_b1_b_85), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_83));
SDFFN u3_mem_reg_b1_b_b0_b (.CK(clk_i), .D(n_8917), .Q(u3_mem_b1_b), .SO(u3_mem_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_85));
SDFFN u8_mem_reg_b1_b_b27_b (.CK(clk_i), .D(n_8914), .Q(u8_mem_b1_b_86), .SO(u8_mem_b1_b_86), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b));
SDFFN u3_mem_reg_b1_b_b10_b (.CK(clk_i), .D(n_8912), .Q(u3_mem_b1_b_69), .SO(u3_mem_b1_b_69), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_86));
SDFFN u8_mem_reg_b1_b_b29_b (.CK(clk_i), .D(n_8910), .Q(u8_mem_b1_b_88), .SO(u8_mem_b1_b_88), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_69));
SDFFN u8_mem_reg_b1_b_b2_b (.CK(clk_i), .D(n_8907), .Q(u8_mem_b1_b_61), .SO(u8_mem_b1_b_61), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_88));
SDFFN u8_mem_reg_b1_b_b30_b (.CK(clk_i), .D(n_8906), .Q(u8_mem_b1_b_89), .SO(u8_mem_b1_b_89), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_61));
SDFFN u8_mem_reg_b1_b_b31_b (.CK(clk_i), .D(n_8351), .Q(u8_mem_b1_b_90), .SO(u8_mem_b1_b_90), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_89));
SDFFN u3_mem_reg_b1_b_b12_b (.CK(clk_i), .D(n_8905), .Q(u3_mem_b1_b_71), .SO(u3_mem_b1_b_71), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_90));
SDFFN u8_mem_reg_b1_b_b4_b (.CK(clk_i), .D(n_8413), .Q(u8_mem_b1_b_63), .SO(u8_mem_b1_b_63), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_71));
SDFFN u3_mem_reg_b1_b_b13_b (.CK(clk_i), .D(n_8901), .Q(u3_mem_b1_b_72), .SO(u3_mem_b1_b_72), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_63));
SDFFN u8_mem_reg_b1_b_b5_b (.CK(clk_i), .D(n_8900), .Q(u8_mem_b1_b_64), .SO(u8_mem_b1_b_64), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_72));
SDFFN u3_mem_reg_b1_b_b14_b (.CK(clk_i), .D(n_9067), .Q(u3_mem_b1_b_73), .SO(u3_mem_b1_b_73), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_64));
SDFFN u8_mem_reg_b1_b_b7_b (.CK(clk_i), .D(n_8899), .Q(u8_mem_b1_b_66), .SO(u8_mem_b1_b_66), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_73));
SDFFN u8_mem_reg_b1_b_b8_b (.CK(clk_i), .D(n_8896), .Q(u8_mem_b1_b_67), .SO(u8_mem_b1_b_67), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_66));
SDFFN u8_mem_reg_b1_b_b9_b (.CK(clk_i), .D(n_8895), .Q(u8_mem_b1_b_68), .SO(u8_mem_b1_b_68), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_67));
SDFFN u8_mem_reg_b2_b_b0_b (.CK(clk_i), .D(n_8892), .Q(u8_mem_b2_b), .SO(u8_mem_b2_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b1_b_68));
SDFFN u3_mem_reg_b1_b_b16_b (.CK(clk_i), .D(n_8893), .Q(u3_mem_b1_b_75), .SO(u3_mem_b1_b_75), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b));
SDFFN u8_mem_reg_b2_b_b10_b (.CK(clk_i), .D(n_8890), .Q(u8_mem_b2_b_38), .SO(u8_mem_b2_b_38), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_75));
SDFFN u8_mem_reg_b2_b_b11_b (.CK(clk_i), .D(n_8886), .Q(u8_mem_b2_b_39), .SO(u8_mem_b2_b_39), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_38));
SDFFN u3_mem_reg_b1_b_b17_b (.CK(clk_i), .D(n_8888), .Q(u3_mem_b1_b_76), .SO(u3_mem_b1_b_76), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_39));
SDFFN u8_mem_reg_b2_b_b12_b (.CK(clk_i), .D(n_8885), .Q(u8_mem_b2_b_40), .SO(u8_mem_b2_b_40), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_76));
SDFFN u3_mem_reg_b1_b_b18_b (.CK(clk_i), .D(n_8883), .Q(u3_mem_b1_b_77), .SO(u3_mem_b1_b_77), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_40));
SDFFN u8_mem_reg_b2_b_b14_b (.CK(clk_i), .D(n_8881), .Q(u8_mem_b2_b_42), .SO(u8_mem_b2_b_42), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_77));
SDFFN u8_mem_reg_b2_b_b15_b (.CK(clk_i), .D(n_8879), .Q(u8_mem_b2_b_43), .SO(u8_mem_b2_b_43), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_42));
SDFFN u8_mem_reg_b2_b_b16_b (.CK(clk_i), .D(n_8878), .Q(u8_mem_b2_b_44), .SO(u8_mem_b2_b_44), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_43));
SDFFN u8_mem_reg_b2_b_b17_b (.CK(clk_i), .D(n_8876), .Q(u8_mem_b2_b_45), .SO(u8_mem_b2_b_45), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_44));
SDFFN u3_mem_reg_b1_b_b1_b (.CK(clk_i), .D(n_8356), .Q(u3_mem_b1_b_60), .SO(u3_mem_b1_b_60), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_45));
SDFFN u8_mem_reg_b2_b_b19_b (.CK(clk_i), .D(n_8872), .Q(u8_mem_b2_b_47), .SO(u8_mem_b2_b_47), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_60));
SDFFN u3_mem_reg_b1_b_b20_b (.CK(clk_i), .D(n_8874), .Q(u3_mem_b1_b_79), .SO(u3_mem_b1_b_79), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_47));
SDFFN u8_mem_reg_b2_b_b1_b (.CK(clk_i), .D(n_8871), .Q(u8_mem_b2_b_29), .SO(u8_mem_b2_b_29), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_79));
SDFFN u3_mem_reg_b1_b_b21_b (.CK(clk_i), .D(n_8870), .Q(u3_mem_b1_b_80), .SO(u3_mem_b1_b_80), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_29));
SDFFN u8_mem_reg_b2_b_b21_b (.CK(clk_i), .D(n_8867), .Q(u8_mem_b2_b_49), .SO(u8_mem_b2_b_49), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_80));
SDFFN u8_mem_reg_b2_b_b22_b (.CK(clk_i), .D(n_8865), .Q(u8_mem_b2_b_50), .SO(u8_mem_b2_b_50), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_49));
SDFFN u8_mem_reg_b2_b_b23_b (.CK(clk_i), .D(n_8864), .Q(u8_mem_b2_b_51), .SO(u8_mem_b2_b_51), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_50));
SDFFN u8_mem_reg_b2_b_b24_b (.CK(clk_i), .D(n_8862), .Q(u8_mem_b2_b_52), .SO(u8_mem_b2_b_52), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_51));
SDFFN u3_mem_reg_b1_b_b23_b (.CK(clk_i), .D(n_9063), .Q(u3_mem_b1_b_82), .SO(u3_mem_b1_b_82), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_52));
SDFFN u8_mem_reg_b2_b_b26_b (.CK(clk_i), .D(n_8859), .Q(u8_mem_b2_b_54), .SO(u8_mem_b2_b_54), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_82));
SDFFN u3_mem_reg_b1_b_b24_b (.CK(clk_i), .D(n_8860), .Q(u3_mem_b1_b_83), .SO(u3_mem_b1_b_83), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_54));
SDFFN u8_mem_reg_b2_b_b27_b (.CK(clk_i), .D(n_8858), .Q(u8_mem_b2_b_55), .SO(u8_mem_b2_b_55), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_83));
SDFFN u3_mem_reg_b1_b_b25_b (.CK(clk_i), .D(n_8857), .Q(u3_mem_b1_b_84), .SO(u3_mem_b1_b_84), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_55));
SDFFN u8_mem_reg_b2_b_b29_b (.CK(clk_i), .D(n_8854), .Q(u8_mem_b2_b_57), .SO(u8_mem_b2_b_57), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_84));
SDFFN u8_mem_reg_b2_b_b2_b (.CK(clk_i), .D(n_8851), .Q(u8_mem_b2_b_30), .SO(u8_mem_b2_b_30), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_57));
SDFFN u8_mem_reg_b2_b_b30_b (.CK(clk_i), .D(n_8850), .Q(u8_mem_b2_b_58), .SO(u8_mem_b2_b_58), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_30));
SDFFN u8_mem_reg_b2_b_b31_b (.CK(clk_i), .D(n_8849), .Q(u8_mem_b2_b_59), .SO(u8_mem_b2_b_59), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_58));
SDFFN u3_mem_reg_b1_b_b27_b (.CK(clk_i), .D(n_8347), .Q(u3_mem_b1_b_86), .SO(u3_mem_b1_b_86), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_59));
SDFFN u4_mem_reg_b0_b_b0_b (.CK(clk_i), .D(n_8837), .Q(u4_mem_b0_b), .SO(u4_mem_b0_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_86));
SDFFN u4_mem_reg_b0_b_b10_b (.CK(clk_i), .D(n_8838), .Q(u4_mem_b0_b_100), .SO(u4_mem_b0_b_100), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b));
SDFFN u4_mem_reg_b0_b_b11_b (.CK(clk_i), .D(n_8836), .Q(u4_mem_b0_b_101), .SO(u4_mem_b0_b_101), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_100));
SDFFN u4_mem_reg_b0_b_b15_b (.CK(clk_i), .D(n_8833), .Q(u4_mem_b0_b_105), .SO(u4_mem_b0_b_105), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_101));
SDFFN u4_mem_reg_b0_b_b18_b (.CK(clk_i), .D(n_8830), .Q(u4_mem_b0_b_108), .SO(u4_mem_b0_b_108), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_105));
SDFFN u4_mem_reg_b0_b_b1_b (.CK(clk_i), .D(n_8829), .Q(u4_mem_b0_b_91), .SO(u4_mem_b0_b_91), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_108));
SDFFN u4_mem_reg_b0_b_b21_b (.CK(clk_i), .D(n_8825), .Q(u4_mem_b0_b_111), .SO(u4_mem_b0_b_111), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_91));
SDFFN u4_mem_reg_b0_b_b25_b (.CK(clk_i), .D(n_8823), .Q(u4_mem_b0_b_115), .SO(u4_mem_b0_b_115), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_111));
SDFFN u4_mem_reg_b0_b_b27_b (.CK(clk_i), .D(n_8821), .Q(u4_mem_b0_b_117), .SO(u4_mem_b0_b_117), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_115));
SDFFN u4_mem_reg_b0_b_b28_b (.CK(clk_i), .D(n_8820), .Q(u4_mem_b0_b_118), .SO(u4_mem_b0_b_118), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_117));
SDFFN u4_mem_reg_b0_b_b26_b (.CK(clk_i), .D(n_8822), .Q(u4_mem_b0_b_116), .SO(u4_mem_b0_b_116), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_118));
SDFFN u4_mem_reg_b0_b_b2_b (.CK(clk_i), .D(n_8817), .Q(u4_mem_b0_b_92), .SO(u4_mem_b0_b_92), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_116));
SDFFN u4_mem_reg_b0_b_b29_b (.CK(clk_i), .D(n_8818), .Q(u4_mem_b0_b_119), .SO(u4_mem_b0_b_119), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_92));
SDFFN u4_mem_reg_b0_b_b3_b (.CK(clk_i), .D(n_8815), .Q(u4_mem_b0_b_93), .SO(u4_mem_b0_b_93), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_119));
SDFFN u4_mem_reg_b0_b_b5_b (.CK(clk_i), .D(n_8813), .Q(u4_mem_b0_b_95), .SO(u4_mem_b0_b_95), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_93));
SDFFN u4_mem_reg_b0_b_b8_b (.CK(clk_i), .D(n_8811), .Q(u4_mem_b0_b_98), .SO(u4_mem_b0_b_98), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_95));
SDFFN u5_mem_reg_b0_b_b10_b (.CK(clk_i), .D(n_8808), .Q(u5_mem_b0_b_100), .SO(u5_mem_b0_b_100), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_98));
SDFFN u5_mem_reg_b0_b_b11_b (.CK(clk_i), .D(n_8807), .Q(u5_mem_b0_b_101), .SO(u5_mem_b0_b_101), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_100));
SDFFN u5_mem_reg_b0_b_b15_b (.CK(clk_i), .D(n_8804), .Q(u5_mem_b0_b_105), .SO(u5_mem_b0_b_105), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_101));
SDFFN u5_mem_reg_b0_b_b18_b (.CK(clk_i), .D(n_8801), .Q(u5_mem_b0_b_108), .SO(u5_mem_b0_b_108), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_105));
SDFFN u5_mem_reg_b0_b_b1_b (.CK(clk_i), .D(n_8800), .Q(u5_mem_b0_b_91), .SO(u5_mem_b0_b_91), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_108));
SDFFN u5_mem_reg_b0_b_b21_b (.CK(clk_i), .D(n_8796), .Q(u5_mem_b0_b_111), .SO(u5_mem_b0_b_111), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_91));
SDFFN u13_intm_r_reg_b8_b (.CK(clk_i), .D(n_8488), .Q(u13_intm_r_b8_b), .SO(u13_intm_r_b8_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_111));
SDFFN u5_mem_reg_b0_b_b26_b (.CK(clk_i), .D(n_8793), .Q(u5_mem_b0_b_116), .SO(u5_mem_b0_b_116), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b8_b));
SDFFN u5_mem_reg_b0_b_b27_b (.CK(clk_i), .D(n_8792), .Q(u5_mem_b0_b_117), .SO(u5_mem_b0_b_117), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_116));
SDFFN u5_mem_reg_b0_b_b25_b (.CK(clk_i), .D(n_8794), .Q(u5_mem_b0_b_115), .SO(u5_mem_b0_b_115), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_117));
SDFFN u5_mem_reg_b0_b_b2_b (.CK(clk_i), .D(n_8788), .Q(u5_mem_b0_b_92), .SO(u5_mem_b0_b_92), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_115));
SDFFN u5_mem_reg_b0_b_b29_b (.CK(clk_i), .D(n_8789), .Q(u5_mem_b0_b_119), .SO(u5_mem_b0_b_119), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_92));
SDFFN u5_mem_reg_b0_b_b3_b (.CK(clk_i), .D(n_8786), .Q(u5_mem_b0_b_93), .SO(u5_mem_b0_b_93), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_119));
SDFFN u5_mem_reg_b0_b_b5_b (.CK(clk_i), .D(n_8784), .Q(u5_mem_b0_b_95), .SO(u5_mem_b0_b_95), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_93));
SDFFN u5_mem_reg_b0_b_b8_b (.CK(clk_i), .D(n_8782), .Q(u5_mem_b0_b_98), .SO(u5_mem_b0_b_98), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_95));
SDFFN u6_mem_reg_b0_b_b10_b (.CK(clk_i), .D(n_8780), .Q(u6_mem_b0_b_100), .SO(u6_mem_b0_b_100), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_98));
SDFFN u6_mem_reg_b0_b_b11_b (.CK(clk_i), .D(n_8779), .Q(u6_mem_b0_b_101), .SO(u6_mem_b0_b_101), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_100));
SDFFN u6_mem_reg_b0_b_b15_b (.CK(clk_i), .D(n_8776), .Q(u6_mem_b0_b_105), .SO(u6_mem_b0_b_105), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_101));
SDFFN u7_mem_reg_b1_b_b21_b (.CK(clk_i), .D(n_9047), .Q(u7_mem_b1_b_80), .SO(u7_mem_b1_b_80), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_105));
SDFFN u6_mem_reg_b0_b_b18_b (.CK(clk_i), .D(n_8773), .Q(u6_mem_b0_b_108), .SO(u6_mem_b0_b_108), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b1_b_80));
SDFFN u6_mem_reg_b0_b_b1_b (.CK(clk_i), .D(n_8772), .Q(u6_mem_b0_b_91), .SO(u6_mem_b0_b_91), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_108));
SDFFN u6_mem_reg_b0_b_b21_b (.CK(clk_i), .D(n_8768), .Q(u6_mem_b0_b_111), .SO(u6_mem_b0_b_111), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_91));
SDFFN u6_mem_reg_b0_b_b26_b (.CK(clk_i), .D(n_8765), .Q(u6_mem_b0_b_116), .SO(u6_mem_b0_b_116), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_111));
SDFFN u6_mem_reg_b0_b_b27_b (.CK(clk_i), .D(n_8764), .Q(u6_mem_b0_b_117), .SO(u6_mem_b0_b_117), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_116));
SDFFN u6_mem_reg_b0_b_b25_b (.CK(clk_i), .D(n_8766), .Q(u6_mem_b0_b_115), .SO(u6_mem_b0_b_115), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_117));
SDFFN u6_mem_reg_b0_b_b2_b (.CK(clk_i), .D(n_8760), .Q(u6_mem_b0_b_92), .SO(u6_mem_b0_b_92), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_115));
SDFFN u6_mem_reg_b0_b_b29_b (.CK(clk_i), .D(n_8761), .Q(u6_mem_b0_b_119), .SO(u6_mem_b0_b_119), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_92));
SDFFN u6_mem_reg_b0_b_b3_b (.CK(clk_i), .D(n_8758), .Q(u6_mem_b0_b_93), .SO(u6_mem_b0_b_93), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_119));
SDFFN u6_mem_reg_b0_b_b5_b (.CK(clk_i), .D(n_8756), .Q(u6_mem_b0_b_95), .SO(u6_mem_b0_b_95), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_93));
SDFFN u6_mem_reg_b0_b_b8_b (.CK(clk_i), .D(n_8754), .Q(u6_mem_b0_b_98), .SO(u6_mem_b0_b_98), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_95));
SDFFN u7_mem_reg_b0_b_b10_b (.CK(clk_i), .D(n_8752), .Q(u7_mem_b0_b_100), .SO(u7_mem_b0_b_100), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b_98));
SDFFN u7_mem_reg_b0_b_b11_b (.CK(clk_i), .D(n_8751), .Q(u7_mem_b0_b_101), .SO(u7_mem_b0_b_101), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_100));
SDFFN u7_mem_reg_b0_b_b15_b (.CK(clk_i), .D(n_8748), .Q(u7_mem_b0_b_105), .SO(u7_mem_b0_b_105), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_101));
SDFFN u7_mem_reg_b0_b_b18_b (.CK(clk_i), .D(n_8745), .Q(u7_mem_b0_b_108), .SO(u7_mem_b0_b_108), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_105));
SDFFN u7_mem_reg_b0_b_b1_b (.CK(clk_i), .D(n_8744), .Q(u7_mem_b0_b_91), .SO(u7_mem_b0_b_91), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_108));
SDFFN u7_mem_reg_b0_b_b21_b (.CK(clk_i), .D(n_8740), .Q(u7_mem_b0_b_111), .SO(u7_mem_b0_b_111), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_91));
SDFFN u7_mem_reg_b0_b_b25_b (.CK(clk_i), .D(n_8738), .Q(u7_mem_b0_b_115), .SO(u7_mem_b0_b_115), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_111));
SDFFN u7_mem_reg_b0_b_b27_b (.CK(clk_i), .D(n_8736), .Q(u7_mem_b0_b_117), .SO(u7_mem_b0_b_117), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_115));
SDFFN u7_mem_reg_b0_b_b28_b (.CK(clk_i), .D(n_8735), .Q(u7_mem_b0_b_118), .SO(u7_mem_b0_b_118), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_117));
SDFFN u7_mem_reg_b0_b_b26_b (.CK(clk_i), .D(n_8737), .Q(u7_mem_b0_b_116), .SO(u7_mem_b0_b_116), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_118));
SDFFN u7_mem_reg_b0_b_b2_b (.CK(clk_i), .D(n_8732), .Q(u7_mem_b0_b_92), .SO(u7_mem_b0_b_92), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_116));
SDFFN u7_mem_reg_b0_b_b29_b (.CK(clk_i), .D(n_8733), .Q(u7_mem_b0_b_119), .SO(u7_mem_b0_b_119), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_92));
SDFFN u7_mem_reg_b0_b_b3_b (.CK(clk_i), .D(n_8730), .Q(u7_mem_b0_b_93), .SO(u7_mem_b0_b_93), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_119));
SDFFN u7_mem_reg_b0_b_b5_b (.CK(clk_i), .D(n_8728), .Q(u7_mem_b0_b_95), .SO(u7_mem_b0_b_95), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_93));
SDFFN u7_mem_reg_b0_b_b8_b (.CK(clk_i), .D(n_8726), .Q(u7_mem_b0_b_98), .SO(u7_mem_b0_b_98), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_95));
SDFFN u3_mem_reg_b0_b_b10_b (.CK(clk_i), .D(n_8725), .Q(u3_mem_b0_b_100), .SO(u3_mem_b0_b_100), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u7_mem_b0_b_98));
SDFFN u8_mem_reg_b0_b_b10_b (.CK(clk_i), .D(n_8721), .Q(u8_mem_b0_b_100), .SO(u8_mem_b0_b_100), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_100));
SDFFN u8_mem_reg_b0_b_b13_b (.CK(clk_i), .D(n_8718), .Q(u8_mem_b0_b_103), .SO(u8_mem_b0_b_103), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_100));
SDFFN u3_mem_reg_b0_b_b18_b (.CK(clk_i), .D(n_8719), .Q(u3_mem_b0_b_108), .SO(u3_mem_b0_b_108), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_103));
SDFFN u8_mem_reg_b0_b_b14_b (.CK(clk_i), .D(n_8717), .Q(u8_mem_b0_b_104), .SO(u8_mem_b0_b_104), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_108));
SDFFN u3_mem_reg_b0_b_b19_b (.CK(clk_i), .D(n_8839), .Q(u3_mem_b0_b_109), .SO(u3_mem_b0_b_109), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_104));
SDFFN u8_mem_reg_b0_b_b18_b (.CK(clk_i), .D(n_8713), .Q(u8_mem_b0_b_108), .SO(u8_mem_b0_b_108), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_109));
SDFFN u8_mem_reg_b0_b_b19_b (.CK(clk_i), .D(n_8709), .Q(u8_mem_b0_b_109), .SO(u8_mem_b0_b_109), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_108));
SDFFN u3_mem_reg_b0_b_b20_b (.CK(clk_i), .D(n_8711), .Q(u3_mem_b0_b_110), .SO(u3_mem_b0_b_110), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_109));
SDFFN u8_mem_reg_b0_b_b20_b (.CK(clk_i), .D(n_8707), .Q(u8_mem_b0_b_110), .SO(u8_mem_b0_b_110), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_110));
SDFFN u8_mem_reg_b0_b_b21_b (.CK(clk_i), .D(n_8705), .Q(u8_mem_b0_b_111), .SO(u8_mem_b0_b_111), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_110));
SDFFN u3_mem_reg_b0_b_b22_b (.CK(clk_i), .D(n_8842), .Q(u3_mem_b0_b_112), .SO(u3_mem_b0_b_112), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_111));
SDFFN u8_mem_reg_b0_b_b23_b (.CK(clk_i), .D(n_8703), .Q(u8_mem_b0_b_113), .SO(u8_mem_b0_b_113), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_112));
SDFFN u8_mem_reg_b0_b_b24_b (.CK(clk_i), .D(n_8699), .Q(u8_mem_b0_b_114), .SO(u8_mem_b0_b_114), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_113));
SDFFN u8_mem_reg_b0_b_b25_b (.CK(clk_i), .D(n_8698), .Q(u8_mem_b0_b_115), .SO(u8_mem_b0_b_115), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_114));
SDFFN u3_mem_reg_b0_b_b24_b (.CK(clk_i), .D(n_8696), .Q(u3_mem_b0_b_114), .SO(u3_mem_b0_b_114), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_115));
SDFFN u3_mem_reg_b0_b_b25_b (.CK(clk_i), .D(n_8694), .Q(u3_mem_b0_b_115), .SO(u3_mem_b0_b_115), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_114));
SDFFN u3_mem_reg_b0_b_b26_b (.CK(clk_i), .D(n_8810), .Q(u3_mem_b0_b_116), .SO(u3_mem_b0_b_116), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_115));
SDFFN u3_mem_reg_b0_b_b28_b (.CK(clk_i), .D(n_8841), .Q(u3_mem_b0_b_118), .SO(u3_mem_b0_b_118), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_116));
SDFFN u8_mem_reg_b0_b_b7_b (.CK(clk_i), .D(n_8688), .Q(u8_mem_b0_b_97), .SO(u8_mem_b0_b_97), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_118));
SDFFN u8_mem_reg_b0_b_b8_b (.CK(clk_i), .D(n_8687), .Q(u8_mem_b0_b_98), .SO(u8_mem_b0_b_98), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_97));
SDFFN u8_mem_reg_b0_b_b6_b (.CK(clk_i), .D(n_8689), .Q(u8_mem_b0_b_96), .SO(u8_mem_b0_b_96), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_98));
SDFFN u8_mem_reg_b0_b_b9_b (.CK(clk_i), .D(n_8686), .Q(u8_mem_b0_b_99), .SO(u8_mem_b0_b_99), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_96));
SDFFN u3_mem_reg_b0_b_b30_b (.CK(clk_i), .D(n_8685), .Q(u3_mem_b0_b_120), .SO(u3_mem_b0_b_120), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_99));
SDFFN u3_mem_reg_b0_b_b3_b (.CK(clk_i), .D(n_8684), .Q(u3_mem_b0_b_93), .SO(u3_mem_b0_b_93), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_120));
SDFFN u3_mem_reg_b0_b_b8_b (.CK(clk_i), .D(n_8681), .Q(u3_mem_b0_b_98), .SO(u3_mem_b0_b_98), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_93));
SDFFN u7_mem_reg_b1_b_b10_b (.CK(clk_i), .D(n_9065), .Q(u7_mem_b1_b_69), .SO(u7_mem_b1_b_69), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_98));
SDFFNSRN u13_crac_dout_r_reg_b7_b (.CK(clk_i), .D(n_8638), .Q(crac_out_852), .SO(crac_out_852), .SE(scan_enable), .SI(u7_mem_b1_b_69));
SDFFN u6_mem_reg_b2_b_b22_b (.CK(clk_i), .D(n_9132), .Q(u6_mem_b2_b_50), .SO(u6_mem_b2_b_50), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_out_852));
SDFFN u6_mem_reg_b0_b_b0_b (.CK(clk_i), .D(n_8781), .Q(u6_mem_b0_b), .SO(u6_mem_b0_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_50));
SDFFN u6_mem_reg_b3_b_b4_b (.CK(clk_i), .D(n_9079), .Q(u6_mem_b3_b_125), .SO(u6_mem_b3_b_125), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b0_b));
SDFFN u13_intm_r_reg_b26_b (.CK(clk_i), .D(n_8500), .Q(u13_intm_r_b26_b), .SO(u13_intm_r_b26_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_125));
SDFFN u6_mem_reg_b3_b_b2_b (.CK(clk_i), .D(n_9084), .Q(u6_mem_b3_b_123), .SO(u6_mem_b3_b_123), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b26_b));
SDFFN u13_occ0_r_reg_b22_b (.CK(clk_i), .D(n_8549), .Q(oc2_cfg_989), .SO(oc2_cfg_989), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_123));
SDFFN u6_mem_reg_b3_b_b26_b (.CK(clk_i), .D(n_9089), .Q(u6_mem_b3_b_147), .SO(u6_mem_b3_b_147), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc2_cfg_989));
SDFFN u6_mem_reg_b3_b_b22_b (.CK(clk_i), .D(n_9094), .Q(u6_mem_b3_b_143), .SO(u6_mem_b3_b_143), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_147));
SDFFN u6_mem_reg_b3_b_b15_b (.CK(clk_i), .D(n_9104), .Q(u6_mem_b3_b_136), .SO(u6_mem_b3_b_136), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_143));
SDFFN u5_mem_reg_b0_b_b6_b (.CK(clk_i), .D(n_8783), .Q(u5_mem_b0_b_96), .SO(u5_mem_b0_b_96), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_136));
SDFFN u6_mem_reg_b3_b_b19_b (.CK(clk_i), .D(n_9099), .Q(u6_mem_b3_b_140), .SO(u6_mem_b3_b_140), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_96));
SDFFN u5_mem_reg_b0_b_b30_b (.CK(clk_i), .D(n_8787), .Q(u5_mem_b0_b_120), .SO(u5_mem_b0_b_120), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_140));
SDFFN u5_mem_reg_b0_b_b23_b (.CK(clk_i), .D(n_8795), .Q(u5_mem_b0_b_113), .SO(u5_mem_b0_b_113), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_120));
SDFFN u13_crac_r_reg_b2_b (.CK(clk_i), .D(n_8634), .Q(crac_out_863), .SO(crac_out_863), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_113));
SDFFN u6_mem_reg_b2_b_b4_b (.CK(clk_i), .D(n_9118), .Q(u6_mem_b2_b_32), .SO(u6_mem_b2_b_32), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_out_863));
SDFFN u6_mem_reg_b3_b_b11_b (.CK(clk_i), .D(n_9109), .Q(u6_mem_b3_b_132), .SO(u6_mem_b3_b_132), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_32));
SDFFN u6_mem_reg_b2_b_b8_b (.CK(clk_i), .D(n_9114), .Q(u6_mem_b2_b_36), .SO(u6_mem_b2_b_36), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b3_b_132));
SDFFN u6_mem_reg_b2_b_b2_b (.CK(clk_i), .D(n_9122), .Q(u6_mem_b2_b_30), .SO(u6_mem_b2_b_30), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_36));
SDFFN u3_mem_reg_b0_b_b9_b (.CK(clk_i), .D(n_8680), .Q(u3_mem_b0_b_99), .SO(u3_mem_b0_b_99), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_30));
SDFFN u13_occ0_r_reg_b26_b (.CK(clk_i), .D(n_8543), .Q(oc3_cfg_995), .SO(oc3_cfg_995), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_99));
SDFFN u5_mem_reg_b0_b_b28_b (.CK(clk_i), .D(n_8791), .Q(u5_mem_b0_b_118), .SO(u5_mem_b0_b_118), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc3_cfg_995));
SDFFN u13_intm_r_reg_b3_b (.CK(clk_i), .D(n_8493), .Q(u13_intm_r_b3_b), .SO(u13_intm_r_b3_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_118));
SDFFN u6_mem_reg_b2_b_b26_b (.CK(clk_i), .D(n_9128), .Q(u6_mem_b2_b_54), .SO(u6_mem_b2_b_54), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_intm_r_b3_b));
SDFFN u3_mem_reg_b0_b_b4_b (.CK(clk_i), .D(n_8682), .Q(u3_mem_b0_b_94), .SO(u3_mem_b0_b_94), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_54));
SDFFN u5_mem_reg_b0_b_b20_b (.CK(clk_i), .D(n_8798), .Q(u5_mem_b0_b_110), .SO(u5_mem_b0_b_110), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_94));
SDFFN u8_mem_reg_b0_b_b31_b (.CK(clk_i), .D(n_8692), .Q(u8_mem_b0_b_121), .SO(u8_mem_b0_b_121), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_110));
SDFFN u6_mem_reg_b2_b_b15_b (.CK(clk_i), .D(n_9142), .Q(u6_mem_b2_b_43), .SO(u6_mem_b2_b_43), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_121));
SDFFN u6_mem_reg_b1_b_b15_b (.CK(clk_i), .D(n_9185), .Q(u6_mem_b1_b_74), .SO(u6_mem_b1_b_74), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_43));
SDFFN u6_mem_reg_b2_b_b19_b (.CK(clk_i), .D(n_9137), .Q(u6_mem_b2_b_47), .SO(u6_mem_b2_b_47), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_74));
SDFFN u6_mem_reg_b2_b_b11_b (.CK(clk_i), .D(n_9147), .Q(u6_mem_b2_b_39), .SO(u6_mem_b2_b_39), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_47));
SDFFN u5_mem_reg_b0_b_b17_b (.CK(clk_i), .D(n_8803), .Q(u5_mem_b0_b_107), .SO(u5_mem_b0_b_107), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b2_b_39));
SDFFN u13_occ0_r_reg_b19_b (.CK(clk_i), .D(n_8556), .Q(oc2_cfg_986), .SO(oc2_cfg_986), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_107));
SDFFN u5_mem_reg_b0_b_b12_b (.CK(clk_i), .D(n_8806), .Q(u5_mem_b0_b_102), .SO(u5_mem_b0_b_102), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc2_cfg_986));
SDFFN u6_mem_reg_b1_b_b26_b (.CK(clk_i), .D(n_9168), .Q(u6_mem_b1_b_85), .SO(u6_mem_b1_b_85), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b_102));
SDFFN u4_mem_reg_b0_b_b6_b (.CK(clk_i), .D(n_8812), .Q(u4_mem_b0_b_96), .SO(u4_mem_b0_b_96), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_85));
SDFFN u6_mem_reg_b1_b_b4_b (.CK(clk_i), .D(n_9156), .Q(u6_mem_b1_b_63), .SO(u6_mem_b1_b_63), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_96));
SDFFN u6_mem_reg_b1_b_b8_b (.CK(clk_i), .D(n_9151), .Q(u6_mem_b1_b_67), .SO(u6_mem_b1_b_67), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_63));
SDFFN u6_mem_reg_b1_b_b2_b (.CK(clk_i), .D(n_9162), .Q(u6_mem_b1_b_61), .SO(u6_mem_b1_b_61), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_67));
SDFFN u5_mem_reg_b0_b_b0_b (.CK(clk_i), .D(n_8809), .Q(u5_mem_b0_b), .SO(u5_mem_b0_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_61));
SDFFN u6_mem_reg_b1_b_b22_b (.CK(clk_i), .D(n_9173), .Q(u6_mem_b1_b_81), .SO(u6_mem_b1_b_81), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b0_b));
SDFFN u8_mem_reg_b0_b_b3_b (.CK(clk_i), .D(n_8691), .Q(u8_mem_b0_b_93), .SO(u8_mem_b0_b_93), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_81));
SDFFN u4_mem_reg_b0_b_b30_b (.CK(clk_i), .D(n_8816), .Q(u4_mem_b0_b_120), .SO(u4_mem_b0_b_120), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_93));
SDFFN u8_mem_reg_b0_b_b16_b (.CK(clk_i), .D(n_8714), .Q(u8_mem_b0_b_106), .SO(u8_mem_b0_b_106), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_120));
SDFFN u5_mem_reg_b3_b_b8_b (.CK(clk_i), .D(n_9199), .Q(u5_mem_b3_b_129), .SO(u5_mem_b3_b_129), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_106));
SDFFN u6_mem_reg_b1_b_b11_b (.CK(clk_i), .D(n_9190), .Q(u6_mem_b1_b_70), .SO(u6_mem_b1_b_70), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_129));
SDFFN u5_mem_reg_b3_b_b4_b (.CK(clk_i), .D(n_9204), .Q(u5_mem_b3_b_125), .SO(u5_mem_b3_b_125), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u6_mem_b1_b_70));
SDFFN u8_mem_reg_b0_b_b2_b (.CK(clk_i), .D(n_8693), .Q(u8_mem_b0_b_92), .SO(u8_mem_b0_b_92), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_125));
SDFFN u5_mem_reg_b2_b_b8_b (.CK(clk_i), .D(n_9239), .Q(u5_mem_b2_b_36), .SO(u5_mem_b2_b_36), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_92));
SDFFN u4_mem_reg_b0_b_b23_b (.CK(clk_i), .D(n_8824), .Q(u4_mem_b0_b_113), .SO(u4_mem_b0_b_113), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_36));
SDFFN u3_mem_reg_b0_b_b23_b (.CK(clk_i), .D(n_8701), .Q(u3_mem_b0_b_113), .SO(u3_mem_b0_b_113), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_113));
SDFFN u4_mem_reg_b0_b_b17_b (.CK(clk_i), .D(n_8832), .Q(u4_mem_b0_b_107), .SO(u4_mem_b0_b_107), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_113));
SDFFN u5_mem_reg_b3_b_b19_b (.CK(clk_i), .D(n_9224), .Q(u5_mem_b3_b_140), .SO(u5_mem_b3_b_140), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_107));
SDFFN u5_mem_reg_b3_b_b26_b (.CK(clk_i), .D(n_9214), .Q(u5_mem_b3_b_147), .SO(u5_mem_b3_b_147), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_140));
SDFFN u5_mem_reg_b3_b_b2_b (.CK(clk_i), .D(n_9209), .Q(u5_mem_b3_b_123), .SO(u5_mem_b3_b_123), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_147));
SDFFN u5_mem_reg_b3_b_b22_b (.CK(clk_i), .D(n_9219), .Q(u5_mem_b3_b_143), .SO(u5_mem_b3_b_143), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_123));
SDFFN u5_mem_reg_b3_b_b15_b (.CK(clk_i), .D(n_9229), .Q(u5_mem_b3_b_136), .SO(u5_mem_b3_b_136), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_143));
SDFFN u8_mem_reg_b0_b_b27_b (.CK(clk_i), .D(n_8695), .Q(u8_mem_b0_b_117), .SO(u8_mem_b0_b_117), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_136));
SDFFN u4_mem_reg_b0_b_b20_b (.CK(clk_i), .D(n_8827), .Q(u4_mem_b0_b_110), .SO(u4_mem_b0_b_110), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_117));
SDFFN u5_mem_reg_b3_b_b11_b (.CK(clk_i), .D(n_9234), .Q(u5_mem_b3_b_132), .SO(u5_mem_b3_b_132), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_110));
SDFFN u5_mem_reg_b2_b_b2_b (.CK(clk_i), .D(n_9247), .Q(u5_mem_b2_b_30), .SO(u5_mem_b2_b_30), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b3_b_132));
SDFFN u4_mem_reg_b0_b_b12_b (.CK(clk_i), .D(n_8835), .Q(u4_mem_b0_b_102), .SO(u4_mem_b0_b_102), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_30));
SDFFN u5_mem_reg_b2_b_b26_b (.CK(clk_i), .D(n_9253), .Q(u5_mem_b2_b_54), .SO(u5_mem_b2_b_54), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u4_mem_b0_b_102));
SDFFN u8_mem_reg_b0_b_b22_b (.CK(clk_i), .D(n_8704), .Q(u8_mem_b0_b_112), .SO(u8_mem_b0_b_112), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_54));
SDFFN u13_occ0_r_reg_b15_b (.CK(clk_i), .D(n_8563), .Q(oc1_cfg_980), .SO(oc1_cfg_980), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_112));
SDFFN u5_mem_reg_b1_b_b2_b (.CK(clk_i), .D(n_9287), .Q(u5_mem_b1_b_61), .SO(u5_mem_b1_b_61), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc1_cfg_980));
SDFFN u5_mem_reg_b2_b_b11_b (.CK(clk_i), .D(n_9272), .Q(u5_mem_b2_b_39), .SO(u5_mem_b2_b_39), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_61));
SDFFN u3_mem_reg_b1_b_b26_b (.CK(clk_i), .D(n_8852), .Q(u3_mem_b1_b_85), .SO(u3_mem_b1_b_85), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_39));
SDFFN u5_mem_reg_b2_b_b19_b (.CK(clk_i), .D(n_9262), .Q(u5_mem_b2_b_47), .SO(u5_mem_b2_b_47), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b1_b_85));
SDFFN u5_mem_reg_b2_b_b22_b (.CK(clk_i), .D(n_9257), .Q(u5_mem_b2_b_50), .SO(u5_mem_b2_b_50), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_47));
SDFFN u5_mem_reg_b2_b_b15_b (.CK(clk_i), .D(n_9267), .Q(u5_mem_b2_b_43), .SO(u5_mem_b2_b_43), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_50));
SDFFN u8_mem_reg_b2_b_b3_b (.CK(clk_i), .D(n_8349), .Q(u8_mem_b2_b_31), .SO(u8_mem_b2_b_31), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b2_b_43));
SDFFN u5_mem_reg_b1_b_b8_b (.CK(clk_i), .D(n_9276), .Q(u5_mem_b1_b_67), .SO(u5_mem_b1_b_67), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b2_b_31));
SDFFN u5_mem_reg_b1_b_b4_b (.CK(clk_i), .D(n_9281), .Q(u5_mem_b1_b_63), .SO(u5_mem_b1_b_63), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_67));
SDFFN u8_mem_reg_b0_b_b1_b (.CK(clk_i), .D(n_8708), .Q(u8_mem_b0_b_91), .SO(u8_mem_b0_b_91), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u5_mem_b1_b_63));
SDFFN u13_occ1_r_reg_b11_b (.CK(clk_i), .D(n_8201), .Q(oc5_cfg_1016), .SO(oc5_cfg_1016), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u8_mem_b0_b_91));
SDFFN u3_mem_reg_b0_b_b0_b (.CK(clk_i), .D(n_8253), .Q(u3_mem_b0_b), .SO(u3_mem_b0_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc5_cfg_1016));
SDFFNSRN u14_u8_en_out_l2_reg (.CK(clk_i), .D(n_9359), .Q(u14_u8_en_out_l2), .SO(u14_u8_en_out_l2), .SE(scan_enable), .SI(u3_mem_b0_b));
SDFFNSRN u12_wb_data_o_reg_b4_b (.CK(clk_i), .D(n_8233), .Q(wb_data_o_b4_b), .SO(wb_data_o_b4_b), .SE(scan_enable), .SI(u14_u8_en_out_l2));
SDFFNSRN u12_wb_data_o_reg_b6_b (.CK(clk_i), .D(n_8231), .Q(wb_data_o_b6_b), .SO(wb_data_o_b6_b), .SE(scan_enable), .SI(wb_data_o_b4_b));
SDFFNSRN u12_wb_data_o_reg_b10_b (.CK(clk_i), .D(n_8244), .Q(wb_data_o_b10_b), .SO(wb_data_o_b10_b), .SE(scan_enable), .SI(wb_data_o_b6_b));
SDFFN u13_occ1_r_reg_b8_b (.CK(clk_i), .D(n_8185), .Q(oc5_cfg), .SO(oc5_cfg), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(wb_data_o_b10_b));
SDFFN u13_occ1_r_reg_b0_b (.CK(clk_i), .D(n_8204), .Q(oc4_cfg), .SO(oc4_cfg), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc5_cfg));
SDFFN u13_occ1_r_reg_b10_b (.CK(clk_i), .D(n_8203), .Q(oc5_cfg_1015), .SO(oc5_cfg_1015), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc4_cfg));
SDFFN u13_occ1_r_reg_b12_b (.CK(clk_i), .D(n_8200), .Q(n_8199), .SO(n_8199), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc5_cfg_1015));
SDFFN u13_occ1_r_reg_b13_b (.CK(clk_i), .D(n_8198), .Q(n_8197), .SO(n_8197), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(n_8199));
SDFFN u13_occ1_r_reg_b14_b (.CK(clk_i), .D(n_8196), .Q(oc5_cfg_1019), .SO(oc5_cfg_1019), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(n_8197));
SDFFN u13_occ1_r_reg_b1_b (.CK(clk_i), .D(n_8194), .Q(oc4_cfg_1004), .SO(oc4_cfg_1004), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc5_cfg_1019));
SDFFN u13_occ1_r_reg_b2_b (.CK(clk_i), .D(n_8193), .Q(oc4_cfg_1005), .SO(oc4_cfg_1005), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc4_cfg_1004));
SDFFN u13_occ1_r_reg_b3_b (.CK(clk_i), .D(n_8192), .Q(oc4_cfg_1006), .SO(oc4_cfg_1006), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc4_cfg_1005));
SDFFN u13_occ1_r_reg_b5_b (.CK(clk_i), .D(n_8189), .Q(n_8188), .SO(n_8188), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc4_cfg_1006));
SDFFN u13_occ1_r_reg_b6_b (.CK(clk_i), .D(n_8187), .Q(oc4_cfg_1009), .SO(oc4_cfg_1009), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(n_8188));
SDFFN u13_occ1_r_reg_b7_b (.CK(clk_i), .D(n_8186), .Q(oc4_cfg_1010), .SO(oc4_cfg_1010), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc4_cfg_1009));
SDFFN u3_mem_reg_b0_b_b14_b (.CK(clk_i), .D(n_8252), .Q(u3_mem_b0_b_104), .SO(u3_mem_b0_b_104), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc4_cfg_1010));
SDFFN u3_mem_reg_b0_b_b7_b (.CK(clk_i), .D(n_8249), .Q(u3_mem_b0_b_97), .SO(u3_mem_b0_b_97), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_104));
SDFFNSRN u14_u6_full_empty_r_reg (.CK(clk_i), .D(n_8215), .Q(u14_u6_full_empty_r), .SO(u14_u6_full_empty_r), .SE(scan_enable), .SI(u3_mem_b0_b_97));
SDFFNSRN u14_u8_full_empty_r_reg (.CK(clk_i), .D(n_8213), .Q(u14_u8_full_empty_r), .SO(u14_u8_full_empty_r), .SE(scan_enable), .SI(u14_u6_full_empty_r));
SDFFNSRN u12_wb_data_o_reg_b0_b (.CK(clk_i), .D(n_8245), .Q(wb_data_o_b0_b), .SO(wb_data_o_b0_b), .SE(scan_enable), .SI(u14_u8_full_empty_r));
SDFFNSRN u12_wb_data_o_reg_b14_b (.CK(clk_i), .D(n_8237), .Q(wb_data_o_b14_b), .SO(wb_data_o_b14_b), .SE(scan_enable), .SI(wb_data_o_b0_b));
SDFFNSRN u12_wb_data_o_reg_b13_b (.CK(clk_i), .D(n_8238), .Q(wb_data_o_b13_b), .SO(wb_data_o_b13_b), .SE(scan_enable), .SI(wb_data_o_b14_b));
SDFFNSRN u12_wb_data_o_reg_b12_b (.CK(clk_i), .D(n_8242), .Q(wb_data_o_b12_b), .SO(wb_data_o_b12_b), .SE(scan_enable), .SI(wb_data_o_b13_b));
SDFFNSRN u12_wb_data_o_reg_b11_b (.CK(clk_i), .D(n_8243), .Q(wb_data_o_b11_b), .SO(wb_data_o_b11_b), .SE(scan_enable), .SI(wb_data_o_b12_b));
SDFFNSRN u12_wb_data_o_reg_b9_b (.CK(clk_i), .D(n_8228), .Q(wb_data_o_b9_b), .SO(wb_data_o_b9_b), .SE(scan_enable), .SI(wb_data_o_b11_b));
SDFFNSRN u12_wb_data_o_reg_b7_b (.CK(clk_i), .D(n_8230), .Q(wb_data_o_b7_b), .SO(wb_data_o_b7_b), .SE(scan_enable), .SI(wb_data_o_b9_b));
SDFFNSRN u12_wb_data_o_reg_b15_b (.CK(clk_i), .D(n_8236), .Q(wb_data_o_b15_b), .SO(wb_data_o_b15_b), .SE(scan_enable), .SI(wb_data_o_b7_b));
SDFFNSRN u12_wb_data_o_reg_b5_b (.CK(clk_i), .D(n_8232), .Q(wb_data_o_b5_b), .SO(wb_data_o_b5_b), .SE(scan_enable), .SI(wb_data_o_b15_b));
SDFFNSRN u12_wb_data_o_reg_b3_b (.CK(clk_i), .D(n_8234), .Q(wb_data_o_b3_b), .SO(wb_data_o_b3_b), .SE(scan_enable), .SI(wb_data_o_b5_b));
SDFFNSRN u12_wb_data_o_reg_b8_b (.CK(clk_i), .D(n_8229), .Q(wb_data_o_b8_b), .SO(wb_data_o_b8_b), .SE(scan_enable), .SI(wb_data_o_b3_b));
SDFFNSRN u12_wb_data_o_reg_b2_b (.CK(clk_i), .D(n_8235), .Q(wb_data_o_b2_b), .SO(wb_data_o_b2_b), .SE(scan_enable), .SI(wb_data_o_b8_b));
SDFFN u13_occ1_r_reg_b9_b (.CK(clk_i), .D(n_8184), .Q(oc5_cfg_1014), .SO(oc5_cfg_1014), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(wb_data_o_b2_b));
SDFFN u13_occ1_r_reg_b15_b (.CK(clk_i), .D(n_8195), .Q(oc5_cfg_1020), .SO(oc5_cfg_1020), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc5_cfg_1014));
SDFFN u3_mem_reg_b0_b_b31_b (.CK(clk_i), .D(n_8250), .Q(u3_mem_b0_b_121), .SO(u3_mem_b0_b_121), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(oc5_cfg_1020));
SDFFN u13_occ1_r_reg_b4_b (.CK(clk_i), .D(n_8191), .Q(n_8190), .SO(n_8190), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u3_mem_b0_b_121));
SDFFNSRN u14_u7_en_out_l2_reg (.CK(clk_i), .D(n_8679), .Q(u14_u7_en_out_l2), .SO(u14_u7_en_out_l2), .SE(scan_enable), .SI(n_8190));
SDFFNSRN u14_u7_full_empty_r_reg (.CK(clk_i), .D(n_7557), .Q(u14_u7_full_empty_r), .SO(u14_u7_full_empty_r), .SE(scan_enable), .SI(u14_u7_en_out_l2));
SDFFNSRN u13_ac97_rst_force_reg (.CK(clk_i), .D(n_7523), .Q(ac97_rst_force), .SO(ac97_rst_force), .SE(scan_enable), .SI(u14_u7_full_empty_r));
SDFFNSRN u13_resume_req_reg (.CK(clk_i), .D(n_7522), .Q(resume_req), .SO(resume_req), .SE(scan_enable), .SI(ac97_rst_force));
SDFFNSRN u14_u6_en_out_l2_reg (.CK(clk_i), .D(n_9352), .Q(u14_u6_en_out_l2), .SO(u14_u6_en_out_l2), .SE(scan_enable), .SI(resume_req));
SDFFNSRN u12_wb_data_o_reg_b31_b (.CK(clk_i), .D(n_7450), .Q(wb_data_o_b31_b), .SO(wb_data_o_b31_b), .SE(scan_enable), .SI(u14_u6_en_out_l2));
SDFFNSRN u12_wb_data_o_reg_b23_b (.CK(clk_i), .D(n_7482), .Q(wb_data_o_b23_b), .SO(wb_data_o_b23_b), .SE(scan_enable), .SI(wb_data_o_b31_b));
SDFFNSRN u12_wb_data_o_reg_b22_b (.CK(clk_i), .D(n_7483), .Q(wb_data_o_b22_b), .SO(wb_data_o_b22_b), .SE(scan_enable), .SI(wb_data_o_b23_b));
SDFFNSRN u12_wb_data_o_reg_b21_b (.CK(clk_i), .D(n_7484), .Q(wb_data_o_b21_b), .SO(wb_data_o_b21_b), .SE(scan_enable), .SI(wb_data_o_b22_b));
SDFFNSRN u12_wb_data_o_reg_b16_b (.CK(clk_i), .D(n_7488), .Q(wb_data_o_b16_b), .SO(wb_data_o_b16_b), .SE(scan_enable), .SI(wb_data_o_b21_b));
SDFFNSRN u12_wb_data_o_reg_b20_b (.CK(clk_i), .D(n_7485), .Q(wb_data_o_b20_b), .SO(wb_data_o_b20_b), .SE(scan_enable), .SI(wb_data_o_b16_b));
SDFFNSRN u12_wb_data_o_reg_b19_b (.CK(clk_i), .D(n_7486), .Q(wb_data_o_b19_b), .SO(wb_data_o_b19_b), .SE(scan_enable), .SI(wb_data_o_b20_b));
SDFFNSRN u12_wb_data_o_reg_b17_b (.CK(clk_i), .D(n_7487), .Q(wb_data_o_b17_b), .SO(wb_data_o_b17_b), .SE(scan_enable), .SI(wb_data_o_b19_b));
SDFFNSRN u12_wb_data_o_reg_b24_b (.CK(clk_i), .D(n_7457), .Q(wb_data_o_b24_b), .SO(wb_data_o_b24_b), .SE(scan_enable), .SI(wb_data_o_b17_b));
SDFFNSRN u12_wb_data_o_reg_b30_b (.CK(clk_i), .D(n_7451), .Q(wb_data_o_b30_b), .SO(wb_data_o_b30_b), .SE(scan_enable), .SI(wb_data_o_b24_b));
SDFFNSRN u12_wb_data_o_reg_b28_b (.CK(clk_i), .D(n_7453), .Q(wb_data_o_b28_b), .SO(wb_data_o_b28_b), .SE(scan_enable), .SI(wb_data_o_b30_b));
SDFFNSRN u12_wb_data_o_reg_b27_b (.CK(clk_i), .D(n_7454), .Q(wb_data_o_b27_b), .SO(wb_data_o_b27_b), .SE(scan_enable), .SI(wb_data_o_b28_b));
SDFFNSRN u12_wb_data_o_reg_b26_b (.CK(clk_i), .D(n_7455), .Q(wb_data_o_b26_b), .SO(wb_data_o_b26_b), .SE(scan_enable), .SI(wb_data_o_b27_b));
SDFFNSRN u12_wb_data_o_reg_b29_b (.CK(clk_i), .D(n_7452), .Q(wb_data_o_b29_b), .SO(wb_data_o_b29_b), .SE(scan_enable), .SI(wb_data_o_b26_b));
SDFFNSRN u12_wb_data_o_reg_b25_b (.CK(clk_i), .D(n_7456), .Q(wb_data_o_b25_b), .SO(wb_data_o_b25_b), .SE(scan_enable), .SI(wb_data_o_b29_b));
SDFFNSRN u12_wb_data_o_reg_b18_b (.CK(clk_i), .D(n_7476), .Q(wb_data_o_b18_b), .SO(wb_data_o_b18_b), .SE(scan_enable), .SI(wb_data_o_b25_b));
SDFFN u4_empty_reg (.CK(clk_i), .D(n_7513), .Q(o4_empty), .SO(o4_empty), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(wb_data_o_b18_b));
SDFFN u6_empty_reg (.CK(clk_i), .D(n_7512), .Q(o7_empty), .SO(o7_empty), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(o4_empty));
SDFFNSRN u15_crac_we_r_reg (.CK(clk_i), .D(n_8643), .Q(u15_crac_we_r), .SO(u15_crac_we_r), .SE(scan_enable), .SI(o7_empty));
SDFFN u3_empty_reg (.CK(clk_i), .D(n_7436), .Q(o3_empty), .SO(o3_empty), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u15_crac_we_r));
SDFFN u5_empty_reg (.CK(clk_i), .D(n_7438), .Q(o6_empty), .SO(o6_empty), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(o3_empty));
SDFFN u7_empty_reg (.CK(clk_i), .D(n_7437), .Q(o8_empty), .SO(o8_empty), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(o6_empty));
SDFFN u8_empty_reg (.CK(clk_i), .D(n_7435), .Q(o9_empty), .SO(o9_empty), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(o8_empty));
SDFFNSRN u10_rp_reg_b2_b (.CK(clk_i), .D(n_7372), .Q(u10_rp_b2_b), .SO(u10_rp_b2_b), .SE(scan_enable), .SI(o9_empty));
SDFFNSRN u11_rp_reg_b2_b (.CK(clk_i), .D(n_7373), .Q(u11_rp_b2_b), .SO(u11_rp_b2_b), .SE(scan_enable), .SI(u10_rp_b2_b));
SDFFN u23_int_set_reg_b1_b (.CK(clk_i), .D(n_7364), .Q(ic0_int_set_719), .SO(ic0_int_set_719), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u11_rp_b2_b));
SDFFN u24_int_set_reg_b1_b (.CK(clk_i), .D(n_7363), .Q(ic1_int_set_721), .SO(ic1_int_set_721), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic0_int_set_719));
SDFFNSRN u11_rp_reg_b1_b (.CK(clk_i), .D(n_7375), .Q(u11_rp_b1_b), .SO(u11_rp_b1_b), .SE(scan_enable), .SI(ic1_int_set_721));
SDFFNSRN u9_rp_reg_b1_b (.CK(clk_i), .D(n_7377), .Q(u9_rp_b1_b), .SO(u9_rp_b1_b), .SE(scan_enable), .SI(u11_rp_b1_b));
SDFFNSRN u10_rp_reg_b1_b (.CK(clk_i), .D(n_7376), .Q(u10_rp_b1_b), .SO(u10_rp_b1_b), .SE(scan_enable), .SI(u9_rp_b1_b));
SDFFNSRN u11_rp_reg_b0_b (.CK(clk_i), .D(n_7371), .Q(u11_rp_b0_b), .SO(u11_rp_b0_b), .SE(scan_enable), .SI(u10_rp_b1_b));
SDFFNSRN u9_rp_reg_b0_b (.CK(clk_i), .D(n_7369), .Q(u9_rp_b0_b), .SO(u9_rp_b0_b), .SE(scan_enable), .SI(u11_rp_b0_b));
SDFFNSRN u9_rp_reg_b2_b (.CK(clk_i), .D(n_7374), .Q(u9_rp_b2_b), .SO(u9_rp_b2_b), .SE(scan_enable), .SI(u9_rp_b0_b));
SDFFNSRN u10_rp_reg_b0_b (.CK(clk_i), .D(n_7366), .Q(u10_rp_b0_b), .SO(u10_rp_b0_b), .SE(scan_enable), .SI(u9_rp_b2_b));
SDFFN u25_int_set_reg_b1_b (.CK(clk_i), .D(n_7280), .Q(ic2_int_set_723), .SO(ic2_int_set_723), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u10_rp_b0_b));
SDFFN valid_s_reg (.CK(clk_i), .D(valid_s1), .Q(valid_s), .SO(valid_s), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(ic2_int_set_723));
SDFFN in_valid_s_reg_b0_b (.CK(clk_i), .D(in_valid_s1), .Q(in_valid_s_b0_b), .SO(in_valid_s_b0_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(valid_s));
SDFFNSRN u12_o7_we_reg (.CK(clk_i), .D(n_7020), .Q(o7_we), .SO(o7_we), .SE(scan_enable), .SI(in_valid_s_b0_b));
SDFFNSRN u12_o3_we_reg (.CK(clk_i), .D(n_7028), .Q(o3_we), .SO(o3_we), .SE(scan_enable), .SI(o7_we));
SDFFNSRN u12_o4_we_reg (.CK(clk_i), .D(n_7027), .Q(o4_we), .SO(o4_we), .SE(scan_enable), .SI(o3_we));
SDFFNSRN u12_o6_we_reg (.CK(clk_i), .D(n_7026), .Q(o6_we), .SO(o6_we), .SE(scan_enable), .SI(o4_we));
SDFFNSRN u12_o8_we_reg (.CK(clk_i), .D(n_7024), .Q(o8_we), .SO(o8_we), .SE(scan_enable), .SI(o6_we));
SDFFNSRN u12_o9_we_reg (.CK(clk_i), .D(n_7023), .Q(o9_we), .SO(o9_we), .SE(scan_enable), .SI(o8_we));
SDFFN in_valid_s_reg_b2_b (.CK(clk_i), .D(in_valid_s_2), .Q(in_valid_s_b2_b), .SO(in_valid_s_b2_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(o9_we));
SDFFN u2_to_cnt_reg_b5_b (.CK(clk_i), .D(n_7033), .Q(u2_to_cnt_b5_b), .SO(u2_to_cnt_b5_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(in_valid_s_b2_b));
SDFFNSRN u13_int_reg (.CK(clk_i), .D(n_7021), .Q(int_o), .SO(int_o), .SE(scan_enable), .SI(u2_to_cnt_b5_b));
SDFFN u13_ints_r_reg_b21_b (.CK(clk_i), .D(n_6753), .Q(u13_ints_r_b21_b), .SO(u13_ints_r_b21_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(int_o));
SDFFN u13_ints_r_reg_b0_b (.CK(clk_i), .D(n_6739), .Q(u13_ints_r_b0_b), .SO(u13_ints_r_b0_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b21_b));
SDFFN u13_ints_r_reg_b27_b (.CK(clk_i), .D(n_6755), .Q(u13_ints_r_b27_b), .SO(u13_ints_r_b27_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b0_b));
SDFFN u13_ints_r_reg_b15_b (.CK(clk_i), .D(n_6744), .Q(u13_ints_r_b15_b), .SO(u13_ints_r_b15_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b27_b));
SDFFN in_valid_s_reg_b1_b (.CK(clk_i), .D(in_valid_s_1), .Q(in_valid_s_b1_b), .SO(in_valid_s_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b15_b));
SDFFNSRN valid_s1_reg (.CK(clk_i), .D(valid), .Q(valid_s1), .SO(valid_s1), .SE(scan_enable), .SI(in_valid_s_b1_b));
SDFFNSRN in_valid_s1_reg_b0_b (.CK(clk_i), .D(in_valid), .Q(in_valid_s1), .SO(in_valid_s1), .SE(scan_enable), .SI(valid_s1));
SDFFN u2_to_cnt_reg_b3_b (.CK(clk_i), .D(n_6065), .Q(u2_to_cnt_b3_b), .SO(u2_to_cnt_b3_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(in_valid_s1));
SDFFNSRN u2_res_cnt_reg_b3_b (.CK(clk_i), .D(n_6067), .Q(u2_res_cnt_b3_b), .SO(u2_res_cnt_b3_b), .SE(scan_enable), .SI(u2_to_cnt_b3_b));
SDFFN u2_to_cnt_reg_b4_b (.CK(clk_i), .D(n_6733), .Q(n_4088), .SO(n_4088), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u2_res_cnt_b3_b));
SDFFNSRN u12_wb_ack_o_reg (.CK(clk_i), .D(n_6716), .Q(wb_ack_o), .SO(wb_ack_o), .SE(scan_enable), .SI(n_4088));
SDFFN u13_ints_r_reg_b10_b (.CK(clk_i), .D(n_6740), .Q(u13_ints_r_b10_b), .SO(u13_ints_r_b10_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(wb_ack_o));
SDFFN u13_ints_r_reg_b12_b (.CK(clk_i), .D(n_6742), .Q(u13_ints_r_b12_b), .SO(u13_ints_r_b12_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b10_b));
SDFFN u13_ints_r_reg_b13_b (.CK(clk_i), .D(n_6741), .Q(u13_ints_r_b13_b), .SO(u13_ints_r_b13_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b12_b));
SDFFN u13_ints_r_reg_b16_b (.CK(clk_i), .D(n_6746), .Q(u13_ints_r_b16_b), .SO(u13_ints_r_b16_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b13_b));
SDFFN u13_ints_r_reg_b18_b (.CK(clk_i), .D(n_6672), .Q(u13_ints_r_b18_b), .SO(u13_ints_r_b18_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b16_b));
SDFFN u13_ints_r_reg_b19_b (.CK(clk_i), .D(n_6747), .Q(u13_ints_r_b19_b), .SO(u13_ints_r_b19_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b18_b));
SDFFN u13_ints_r_reg_b22_b (.CK(clk_i), .D(n_6749), .Q(u13_ints_r_b22_b), .SO(u13_ints_r_b22_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b19_b));
SDFFN u13_ints_r_reg_b24_b (.CK(clk_i), .D(n_6751), .Q(u13_ints_r_b24_b), .SO(u13_ints_r_b24_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b22_b));
SDFFN u13_ints_r_reg_b25_b (.CK(clk_i), .D(n_6754), .Q(u13_ints_r_b25_b), .SO(u13_ints_r_b25_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b24_b));
SDFFN u13_ints_r_reg_b28_b (.CK(clk_i), .D(n_6758), .Q(u13_ints_r_b28_b), .SO(u13_ints_r_b28_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b25_b));
SDFFN u13_ints_r_reg_b3_b (.CK(clk_i), .D(n_6759), .Q(u13_ints_r_b3_b), .SO(u13_ints_r_b3_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b28_b));
SDFFN u13_ints_r_reg_b4_b (.CK(clk_i), .D(n_6671), .Q(u13_ints_r_b4_b), .SO(u13_ints_r_b4_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b3_b));
SDFFN u13_ints_r_reg_b7_b (.CK(clk_i), .D(n_6063), .Q(u13_ints_r_b7_b), .SO(u13_ints_r_b7_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b4_b));
SDFFN u13_ints_r_reg_b6_b (.CK(clk_i), .D(n_6062), .Q(u13_ints_r_b6_b), .SO(u13_ints_r_b6_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b7_b));
SDFFN u13_ints_r_reg_b9_b (.CK(clk_i), .D(n_6064), .Q(u13_ints_r_b9_b), .SO(u13_ints_r_b9_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b6_b));
SDFFN u2_to_cnt_reg_b2_b (.CK(clk_i), .D(n_6054), .Q(n_1819), .SO(n_1819), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u13_ints_r_b9_b));
SDFFNSRN u4_status_reg_b1_b (.CK(clk_i), .D(n_6050), .Q(o4_status_972), .SO(o4_status_972), .SE(scan_enable), .SI(n_1819));
SDFFNSRN u5_status_reg_b1_b (.CK(clk_i), .D(n_6048), .Q(o6_status_982), .SO(o6_status_982), .SE(scan_enable), .SI(o4_status_972));
SDFFNSRN u12_rf_we_reg (.CK(clk_i), .D(n_6041), .Q(rf_we), .SO(rf_we), .SE(scan_enable), .SI(o6_status_982));
SDFFNSRN u2_res_cnt_reg_b0_b (.CK(clk_i), .D(n_6053), .Q(u2_res_cnt_b0_b), .SO(u2_res_cnt_b0_b), .SE(scan_enable), .SI(rf_we));
SDFFNSRN in_valid_s1_reg_b2_b (.CK(clk_i), .D(in_valid_9), .Q(in_valid_s_2), .SO(in_valid_s_2), .SE(scan_enable), .SI(u2_res_cnt_b0_b));
SDFFN u2_to_cnt_reg_b0_b (.CK(clk_i), .D(n_5976), .Q(u2_to_cnt_b0_b), .SO(u2_to_cnt_b0_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(in_valid_s_2));
SDFFN u2_to_cnt_reg_b1_b (.CK(clk_i), .D(n_6025), .Q(u2_to_cnt_b1_b), .SO(u2_to_cnt_b1_b), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(u2_to_cnt_b0_b));
SDFFNSRN u2_res_cnt_reg_b2_b (.CK(clk_i), .D(n_5628), .Q(u2_res_cnt_b2_b), .SO(u2_res_cnt_b2_b), .SE(scan_enable), .SI(u2_to_cnt_b1_b));
SDFFNSRN u2_res_cnt_reg_b1_b (.CK(clk_i), .D(n_5627), .Q(u2_res_cnt_b1_b), .SO(u2_res_cnt_b1_b), .SE(scan_enable), .SI(u2_res_cnt_b2_b));
SDFFNSRN u3_status_reg_b1_b (.CK(clk_i), .D(n_5621), .Q(o3_status_962), .SO(o3_status_962), .SE(scan_enable), .SI(u2_res_cnt_b1_b));
SDFFNSRN u6_status_reg_b1_b (.CK(clk_i), .D(n_5619), .Q(o7_status_992), .SO(o7_status_992), .SE(scan_enable), .SI(o3_status_962));
SDFFNSRN u7_status_reg_b1_b (.CK(clk_i), .D(n_5617), .Q(o8_status_1002), .SO(o8_status_1002), .SE(scan_enable), .SI(o7_status_992));
SDFFNSRN u8_status_reg_b1_b (.CK(clk_i), .D(n_5623), .Q(o9_status_1012), .SO(o9_status_1012), .SE(scan_enable), .SI(o8_status_1002));
SDFFNSRN u11_status_reg_b1_b (.CK(clk_i), .D(n_5638), .Q(i6_status_1042), .SO(i6_status_1042), .SE(scan_enable), .SI(o9_status_1012));
SDFFNSRN u10_empty_reg (.CK(clk_i), .D(n_5612), .Q(i4_empty), .SO(i4_empty), .SE(scan_enable), .SI(i6_status_1042));
SDFFNSRN u9_empty_reg (.CK(clk_i), .D(n_5613), .Q(i3_empty), .SO(i3_empty), .SE(scan_enable), .SI(i4_empty));
SDFFNSRN in_valid_s1_reg_b1_b (.CK(clk_i), .D(in_valid_8), .Q(in_valid_s_1), .SO(in_valid_s_1), .SE(scan_enable), .SI(i3_empty));
SDFFNSRN u12_we1_reg (.CK(clk_i), .D(n_5361), .Q(u12_we1), .SO(u12_we1), .SE(scan_enable), .SI(in_valid_s_1));
SDFFNSRN u10_status_reg_b1_b (.CK(clk_i), .D(n_5431), .Q(i4_status_1032), .SO(i4_status_1032), .SE(scan_enable), .SI(u12_we1));
SDFFNSRN u9_status_reg_b1_b (.CK(clk_i), .D(n_5449), .Q(i3_status_1022), .SO(i3_status_1022), .SE(scan_enable), .SI(i4_status_1032));
SDFFNSRN u11_empty_reg (.CK(clk_i), .D(n_5383), .Q(i6_empty), .SO(i6_empty), .SE(scan_enable), .SI(i3_status_1022));
SDFFN u11_full_reg (.CK(clk_i), .D(n_5443), .Q(i6_full), .SO(i6_full), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(i6_empty));
SDFFNSRN u10_dout_reg_b14_b (.CK(clk_i), .D(n_5382), .Q(i4_dout_608), .SO(i4_dout_608), .SE(scan_enable), .SI(i6_full));
SDFFNSRN u10_dout_reg_b15_b (.CK(clk_i), .D(n_5393), .Q(i4_dout_609), .SO(i4_dout_609), .SE(scan_enable), .SI(i4_dout_608));
SDFFNSRN u10_dout_reg_b17_b (.CK(clk_i), .D(n_5392), .Q(i4_dout_611), .SO(i4_dout_611), .SE(scan_enable), .SI(i4_dout_609));
SDFFNSRN u10_dout_reg_b18_b (.CK(clk_i), .D(n_5391), .Q(i4_dout_612), .SO(i4_dout_612), .SE(scan_enable), .SI(i4_dout_611));
SDFFNSRN u10_dout_reg_b19_b (.CK(clk_i), .D(n_5390), .Q(i4_dout_613), .SO(i4_dout_613), .SE(scan_enable), .SI(i4_dout_612));
SDFFNSRN u10_dout_reg_b1_b (.CK(clk_i), .D(n_5389), .Q(i4_dout_595), .SO(i4_dout_595), .SE(scan_enable), .SI(i4_dout_613));
SDFFNSRN u10_dout_reg_b20_b (.CK(clk_i), .D(n_5388), .Q(i4_dout_614), .SO(i4_dout_614), .SE(scan_enable), .SI(i4_dout_595));
SDFFNSRN u10_dout_reg_b21_b (.CK(clk_i), .D(n_5387), .Q(i4_dout_615), .SO(i4_dout_615), .SE(scan_enable), .SI(i4_dout_614));
SDFFNSRN u10_dout_reg_b22_b (.CK(clk_i), .D(n_5386), .Q(i4_dout_616), .SO(i4_dout_616), .SE(scan_enable), .SI(i4_dout_615));
SDFFNSRN u10_dout_reg_b23_b (.CK(clk_i), .D(n_5385), .Q(i4_dout_617), .SO(i4_dout_617), .SE(scan_enable), .SI(i4_dout_616));
SDFFNSRN u12_i4_re_reg (.CK(clk_i), .D(n_4838), .Q(i4_re), .SO(i4_re), .SE(scan_enable), .SI(i4_dout_617));
SDFFN u9_full_reg (.CK(clk_i), .D(n_4852), .Q(i3_full), .SO(i3_full), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(i4_re));
SDFFN u12_i6_re_reg (.CK(clk_i), .D(n_4828), .Q(i6_re), .SO(i6_re), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(i3_full));
SDFFN u12_i3_re_reg (.CK(clk_i), .D(n_4839), .Q(i3_re), .SO(i3_re), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(i6_re));
SDFFNSRN u10_dout_reg_b11_b (.CK(clk_i), .D(n_4823), .Q(i4_dout_605), .SO(i4_dout_605), .SE(scan_enable), .SI(i3_re));
SDFFNSRN u10_dout_reg_b0_b (.CK(clk_i), .D(n_4824), .Q(i4_dout), .SO(i4_dout), .SE(scan_enable), .SI(i4_dout_605));
SDFFNSRN u10_dout_reg_b10_b (.CK(clk_i), .D(n_4807), .Q(i4_dout_604), .SO(i4_dout_604), .SE(scan_enable), .SI(i4_dout));
SDFFNSRN u10_dout_reg_b12_b (.CK(clk_i), .D(n_4822), .Q(i4_dout_606), .SO(i4_dout_606), .SE(scan_enable), .SI(i4_dout_604));
SDFFNSRN u10_dout_reg_b13_b (.CK(clk_i), .D(n_4821), .Q(i4_dout_607), .SO(i4_dout_607), .SE(scan_enable), .SI(i4_dout_606));
SDFFNSRN u10_dout_reg_b25_b (.CK(clk_i), .D(n_4818), .Q(i4_dout_619), .SO(i4_dout_619), .SE(scan_enable), .SI(i4_dout_607));
SDFFNSRN u10_dout_reg_b27_b (.CK(clk_i), .D(n_4817), .Q(i4_dout_621), .SO(i4_dout_621), .SE(scan_enable), .SI(i4_dout_619));
SDFFNSRN u10_dout_reg_b28_b (.CK(clk_i), .D(n_4816), .Q(i4_dout_622), .SO(i4_dout_622), .SE(scan_enable), .SI(i4_dout_621));
SDFFNSRN u10_dout_reg_b29_b (.CK(clk_i), .D(n_4815), .Q(i4_dout_623), .SO(i4_dout_623), .SE(scan_enable), .SI(i4_dout_622));
SDFFNSRN u10_dout_reg_b2_b (.CK(clk_i), .D(n_4806), .Q(i4_dout_596), .SO(i4_dout_596), .SE(scan_enable), .SI(i4_dout_623));
SDFFNSRN u10_dout_reg_b30_b (.CK(clk_i), .D(n_4814), .Q(i4_dout_624), .SO(i4_dout_624), .SE(scan_enable), .SI(i4_dout_596));
SDFFNSRN u10_dout_reg_b3_b (.CK(clk_i), .D(n_4813), .Q(i4_dout_597), .SO(i4_dout_597), .SE(scan_enable), .SI(i4_dout_624));
SDFFNSRN u10_dout_reg_b4_b (.CK(clk_i), .D(n_4812), .Q(i4_dout_598), .SO(i4_dout_598), .SE(scan_enable), .SI(i4_dout_597));
SDFFNSRN u10_dout_reg_b6_b (.CK(clk_i), .D(n_4811), .Q(i4_dout_600), .SO(i4_dout_600), .SE(scan_enable), .SI(i4_dout_598));
SDFFNSRN u10_dout_reg_b7_b (.CK(clk_i), .D(n_4810), .Q(i4_dout_601), .SO(i4_dout_601), .SE(scan_enable), .SI(i4_dout_600));
SDFFNSRN u10_dout_reg_b8_b (.CK(clk_i), .D(n_4809), .Q(i4_dout_602), .SO(i4_dout_602), .SE(scan_enable), .SI(i4_dout_601));
SDFFNSRN u10_dout_reg_b9_b (.CK(clk_i), .D(n_4808), .Q(i4_dout_603), .SO(i4_dout_603), .SE(scan_enable), .SI(i4_dout_602));
SDFFN u10_full_reg (.CK(clk_i), .D(n_4105), .Q(i4_full), .SO(i4_full), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(i4_dout_603));
SDFFNSRN u9_dout_reg_b11_b (.CK(clk_i), .D(n_4065), .Q(i3_dout_574), .SO(i3_dout_574), .SE(scan_enable), .SI(i4_full));
SDFFNSRN u9_dout_reg_b14_b (.CK(clk_i), .D(n_4062), .Q(i3_dout_577), .SO(i3_dout_577), .SE(scan_enable), .SI(i3_dout_574));
SDFFNSRN u9_dout_reg_b18_b (.CK(clk_i), .D(n_4058), .Q(i3_dout_581), .SO(i3_dout_581), .SE(scan_enable), .SI(i3_dout_577));
SDFFNSRN u9_dout_reg_b19_b (.CK(clk_i), .D(n_4057), .Q(i3_dout_582), .SO(i3_dout_582), .SE(scan_enable), .SI(i3_dout_581));
SDFFNSRN u9_dout_reg_b20_b (.CK(clk_i), .D(n_4055), .Q(i3_dout_583), .SO(i3_dout_583), .SE(scan_enable), .SI(i3_dout_582));
SDFFNSRN u9_dout_reg_b21_b (.CK(clk_i), .D(n_4054), .Q(i3_dout_584), .SO(i3_dout_584), .SE(scan_enable), .SI(i3_dout_583));
SDFFNSRN u9_dout_reg_b22_b (.CK(clk_i), .D(n_4053), .Q(i3_dout_585), .SO(i3_dout_585), .SE(scan_enable), .SI(i3_dout_584));
SDFFNSRN u9_dout_reg_b23_b (.CK(clk_i), .D(n_4052), .Q(i3_dout_586), .SO(i3_dout_586), .SE(scan_enable), .SI(i3_dout_585));
SDFFNSRN u9_dout_reg_b24_b (.CK(clk_i), .D(n_4051), .Q(i3_dout_587), .SO(i3_dout_587), .SE(scan_enable), .SI(i3_dout_586));
SDFFNSRN u9_dout_reg_b25_b (.CK(clk_i), .D(n_4039), .Q(i3_dout_588), .SO(i3_dout_588), .SE(scan_enable), .SI(i3_dout_587));
SDFFNSRN u9_dout_reg_b16_b (.CK(clk_i), .D(n_4060), .Q(i3_dout_579), .SO(i3_dout_579), .SE(scan_enable), .SI(i3_dout_588));
SDFFNSRN u10_dout_reg_b16_b (.CK(clk_i), .D(n_4342), .Q(i4_dout_610), .SO(i4_dout_610), .SE(scan_enable), .SI(i3_dout_579));
SDFFNSRN u9_dout_reg_b26_b (.CK(clk_i), .D(n_4050), .Q(i3_dout_589), .SO(i3_dout_589), .SE(scan_enable), .SI(i4_dout_610));
SDFFNSRN u9_dout_reg_b27_b (.CK(clk_i), .D(n_4049), .Q(i3_dout_590), .SO(i3_dout_590), .SE(scan_enable), .SI(i3_dout_589));
SDFFNSRN u9_dout_reg_b28_b (.CK(clk_i), .D(n_4048), .Q(i3_dout_591), .SO(i3_dout_591), .SE(scan_enable), .SI(i3_dout_590));
SDFFNSRN u9_dout_reg_b29_b (.CK(clk_i), .D(n_4047), .Q(i3_dout_592), .SO(i3_dout_592), .SE(scan_enable), .SI(i3_dout_591));
SDFFNSRN u9_dout_reg_b2_b (.CK(clk_i), .D(n_4046), .Q(i3_dout_565), .SO(i3_dout_565), .SE(scan_enable), .SI(i3_dout_592));
SDFFNSRN u9_dout_reg_b30_b (.CK(clk_i), .D(n_4045), .Q(i3_dout_593), .SO(i3_dout_593), .SE(scan_enable), .SI(i3_dout_565));
SDFFNSRN u9_dout_reg_b31_b (.CK(clk_i), .D(n_4044), .Q(i3_dout_594), .SO(i3_dout_594), .SE(scan_enable), .SI(i3_dout_593));
SDFFNSRN u9_dout_reg_b3_b (.CK(clk_i), .D(n_4043), .Q(i3_dout_566), .SO(i3_dout_566), .SE(scan_enable), .SI(i3_dout_594));
SDFFNSRN u9_dout_reg_b4_b (.CK(clk_i), .D(n_4033), .Q(i3_dout_567), .SO(i3_dout_567), .SE(scan_enable), .SI(i3_dout_566));
SDFFNSRN u9_dout_reg_b5_b (.CK(clk_i), .D(n_4042), .Q(i3_dout_568), .SO(i3_dout_568), .SE(scan_enable), .SI(i3_dout_567));
SDFFNSRN u9_dout_reg_b6_b (.CK(clk_i), .D(n_4041), .Q(i3_dout_569), .SO(i3_dout_569), .SE(scan_enable), .SI(i3_dout_568));
SDFFNSRN u9_dout_reg_b7_b (.CK(clk_i), .D(n_4040), .Q(i3_dout_570), .SO(i3_dout_570), .SE(scan_enable), .SI(i3_dout_569));
SDFFNSRN u9_dout_reg_b8_b (.CK(clk_i), .D(n_3999), .Q(i3_dout_571), .SO(i3_dout_571), .SE(scan_enable), .SI(i3_dout_570));
SDFFNSRN u9_dout_reg_b9_b (.CK(clk_i), .D(n_3997), .Q(i3_dout_572), .SO(i3_dout_572), .SE(scan_enable), .SI(i3_dout_571));
SDFFNSRN u10_dout_reg_b24_b (.CK(clk_i), .D(n_4037), .Q(i4_dout_618), .SO(i4_dout_618), .SE(scan_enable), .SI(i3_dout_572));
SDFFNSRN u10_dout_reg_b26_b (.CK(clk_i), .D(n_4034), .Q(i4_dout_620), .SO(i4_dout_620), .SE(scan_enable), .SI(i4_dout_618));
SDFFNSRN u9_dout_reg_b13_b (.CK(clk_i), .D(n_4063), .Q(i3_dout_576), .SO(i3_dout_576), .SE(scan_enable), .SI(i4_dout_620));
SDFFNSRN u11_dout_reg_b0_b (.CK(clk_i), .D(n_4032), .Q(i6_dout), .SO(i6_dout), .SE(scan_enable), .SI(i3_dout_576));
SDFFNSRN u11_dout_reg_b10_b (.CK(clk_i), .D(n_4031), .Q(i6_dout_635), .SO(i6_dout_635), .SE(scan_enable), .SI(i6_dout));
SDFFNSRN u11_dout_reg_b11_b (.CK(clk_i), .D(n_4030), .Q(i6_dout_636), .SO(i6_dout_636), .SE(scan_enable), .SI(i6_dout_635));
SDFFNSRN u11_dout_reg_b12_b (.CK(clk_i), .D(n_4029), .Q(i6_dout_637), .SO(i6_dout_637), .SE(scan_enable), .SI(i6_dout_636));
SDFFNSRN u11_dout_reg_b13_b (.CK(clk_i), .D(n_4028), .Q(i6_dout_638), .SO(i6_dout_638), .SE(scan_enable), .SI(i6_dout_637));
SDFFNSRN u10_dout_reg_b31_b (.CK(clk_i), .D(n_3998), .Q(i4_dout_625), .SO(i4_dout_625), .SE(scan_enable), .SI(i6_dout_638));
SDFFNSRN u11_dout_reg_b14_b (.CK(clk_i), .D(n_4027), .Q(i6_dout_639), .SO(i6_dout_639), .SE(scan_enable), .SI(i4_dout_625));
SDFFNSRN u11_dout_reg_b15_b (.CK(clk_i), .D(n_4026), .Q(i6_dout_640), .SO(i6_dout_640), .SE(scan_enable), .SI(i6_dout_639));
SDFFNSRN u11_dout_reg_b16_b (.CK(clk_i), .D(n_4025), .Q(i6_dout_641), .SO(i6_dout_641), .SE(scan_enable), .SI(i6_dout_640));
SDFFNSRN u11_dout_reg_b17_b (.CK(clk_i), .D(n_4024), .Q(i6_dout_642), .SO(i6_dout_642), .SE(scan_enable), .SI(i6_dout_641));
SDFFNSRN u11_dout_reg_b18_b (.CK(clk_i), .D(n_4023), .Q(i6_dout_643), .SO(i6_dout_643), .SE(scan_enable), .SI(i6_dout_642));
SDFFNSRN u11_dout_reg_b19_b (.CK(clk_i), .D(n_4021), .Q(i6_dout_644), .SO(i6_dout_644), .SE(scan_enable), .SI(i6_dout_643));
SDFFNSRN u10_dout_reg_b5_b (.CK(clk_i), .D(n_4022), .Q(i4_dout_599), .SO(i4_dout_599), .SE(scan_enable), .SI(i6_dout_644));
SDFFNSRN u11_dout_reg_b1_b (.CK(clk_i), .D(n_4020), .Q(i6_dout_626), .SO(i6_dout_626), .SE(scan_enable), .SI(i4_dout_599));
SDFFNSRN u11_dout_reg_b20_b (.CK(clk_i), .D(n_4019), .Q(i6_dout_645), .SO(i6_dout_645), .SE(scan_enable), .SI(i6_dout_626));
SDFFNSRN u11_dout_reg_b21_b (.CK(clk_i), .D(n_4018), .Q(i6_dout_646), .SO(i6_dout_646), .SE(scan_enable), .SI(i6_dout_645));
SDFFNSRN u11_dout_reg_b22_b (.CK(clk_i), .D(n_4017), .Q(i6_dout_647), .SO(i6_dout_647), .SE(scan_enable), .SI(i6_dout_646));
SDFFNSRN u11_dout_reg_b23_b (.CK(clk_i), .D(n_4016), .Q(i6_dout_648), .SO(i6_dout_648), .SE(scan_enable), .SI(i6_dout_647));
SDFFNSRN u11_dout_reg_b24_b (.CK(clk_i), .D(n_4015), .Q(i6_dout_649), .SO(i6_dout_649), .SE(scan_enable), .SI(i6_dout_648));
SDFFNSRN u11_dout_reg_b25_b (.CK(clk_i), .D(n_4014), .Q(i6_dout_650), .SO(i6_dout_650), .SE(scan_enable), .SI(i6_dout_649));
SDFFNSRN u11_dout_reg_b26_b (.CK(clk_i), .D(n_4013), .Q(i6_dout_651), .SO(i6_dout_651), .SE(scan_enable), .SI(i6_dout_650));
SDFFNSRN u11_dout_reg_b27_b (.CK(clk_i), .D(n_4012), .Q(i6_dout_652), .SO(i6_dout_652), .SE(scan_enable), .SI(i6_dout_651));
SDFFNSRN u11_dout_reg_b28_b (.CK(clk_i), .D(n_4011), .Q(i6_dout_653), .SO(i6_dout_653), .SE(scan_enable), .SI(i6_dout_652));
SDFFNSRN u11_dout_reg_b29_b (.CK(clk_i), .D(n_4010), .Q(i6_dout_654), .SO(i6_dout_654), .SE(scan_enable), .SI(i6_dout_653));
SDFFNSRN u11_dout_reg_b2_b (.CK(clk_i), .D(n_4009), .Q(i6_dout_627), .SO(i6_dout_627), .SE(scan_enable), .SI(i6_dout_654));
SDFFNSRN u11_dout_reg_b30_b (.CK(clk_i), .D(n_4008), .Q(i6_dout_655), .SO(i6_dout_655), .SE(scan_enable), .SI(i6_dout_627));
SDFFNSRN u11_dout_reg_b31_b (.CK(clk_i), .D(n_4007), .Q(i6_dout_656), .SO(i6_dout_656), .SE(scan_enable), .SI(i6_dout_655));
SDFFNSRN u11_dout_reg_b3_b (.CK(clk_i), .D(n_4006), .Q(i6_dout_628), .SO(i6_dout_628), .SE(scan_enable), .SI(i6_dout_656));
SDFFNSRN u11_dout_reg_b4_b (.CK(clk_i), .D(n_4005), .Q(i6_dout_629), .SO(i6_dout_629), .SE(scan_enable), .SI(i6_dout_628));
SDFFNSRN u11_dout_reg_b5_b (.CK(clk_i), .D(n_4004), .Q(i6_dout_630), .SO(i6_dout_630), .SE(scan_enable), .SI(i6_dout_629));
SDFFNSRN u11_dout_reg_b6_b (.CK(clk_i), .D(n_4038), .Q(i6_dout_631), .SO(i6_dout_631), .SE(scan_enable), .SI(i6_dout_630));
SDFFNSRN u11_dout_reg_b7_b (.CK(clk_i), .D(n_4003), .Q(i6_dout_632), .SO(i6_dout_632), .SE(scan_enable), .SI(i6_dout_631));
SDFFNSRN u11_dout_reg_b8_b (.CK(clk_i), .D(n_4002), .Q(i6_dout_633), .SO(i6_dout_633), .SE(scan_enable), .SI(i6_dout_632));
SDFFNSRN u11_dout_reg_b9_b (.CK(clk_i), .D(n_4001), .Q(i6_dout_634), .SO(i6_dout_634), .SE(scan_enable), .SI(i6_dout_633));
SDFFNSRN u9_dout_reg_b15_b (.CK(clk_i), .D(n_4061), .Q(i3_dout_578), .SO(i3_dout_578), .SE(scan_enable), .SI(i6_dout_634));
SDFFNSRN u9_dout_reg_b17_b (.CK(clk_i), .D(n_4059), .Q(i3_dout_580), .SO(i3_dout_580), .SE(scan_enable), .SI(i3_dout_578));
SDFFNSRN u9_dout_reg_b0_b (.CK(clk_i), .D(n_4067), .Q(i3_dout), .SO(i3_dout), .SE(scan_enable), .SI(i3_dout_580));
SDFFNSRN u9_dout_reg_b12_b (.CK(clk_i), .D(n_4064), .Q(i3_dout_575), .SO(i3_dout_575), .SE(scan_enable), .SI(i3_dout));
SDFFNSRN u9_dout_reg_b10_b (.CK(clk_i), .D(n_4066), .Q(i3_dout_573), .SO(i3_dout_573), .SE(scan_enable), .SI(i3_dout_575));
SDFFNSRN u9_dout_reg_b1_b (.CK(clk_i), .D(n_4056), .Q(i3_dout_564), .SO(i3_dout_564), .SE(scan_enable), .SI(i3_dout_573));
SDFFN u12_re2_reg (.CK(clk_i), .D(n_4086), .Q(u12_re2), .SO(u12_re2), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(i3_dout_564));
SDFFNSRN u12_re1_reg (.CK(clk_i), .D(n_2600), .Q(u12_re1), .SO(u12_re1), .SE(scan_enable), .SI(u12_re2));
SDFFNSRN u2_bit_clk_e_reg (.CK(clk_i), .D(n_2589), .Q(u2_bit_clk_e), .SO(u2_bit_clk_e), .SE(scan_enable), .SI(u12_re1));
SDFFNSRN u2_suspended_reg (.CK(clk_i), .D(n_5630), .Q(suspended_o), .SO(suspended_o), .SE(scan_enable), .SI(u2_bit_clk_e));
SDFFNSRN u10_status_reg_b0_b (.CK(clk_i), .D(n_3561), .Q(i4_status), .SO(i4_status), .SE(scan_enable), .SI(suspended_o));
SDFFNSRN u9_status_reg_b0_b (.CK(clk_i), .D(n_3563), .Q(i3_status), .SO(i3_status), .SE(scan_enable), .SI(i4_status));
SDFFNSRN u11_status_reg_b0_b (.CK(clk_i), .D(n_1804), .Q(i6_status), .SO(i6_status), .SE(scan_enable), .SI(i3_status));
SDFFNSRN u6_status_reg_b0_b (.CK(clk_i), .D(n_5618), .Q(o7_status), .SO(o7_status), .SE(scan_enable), .SI(i6_status));
SDFFNSRN u3_status_reg_b0_b (.CK(clk_i), .D(n_5620), .Q(o3_status), .SO(o3_status), .SE(scan_enable), .SI(o7_status));
SDFFNSRN u4_status_reg_b0_b (.CK(clk_i), .D(n_6049), .Q(o4_status), .SO(o4_status), .SE(scan_enable), .SI(o3_status));
SDFFNSRN u7_status_reg_b0_b (.CK(clk_i), .D(n_5616), .Q(o8_status), .SO(o8_status), .SE(scan_enable), .SI(o4_status));
SDFFN u15_crac_din_reg_b6_b (.CK(clk_i), .D(n_1196), .Q(crac_din_697), .SO(crac_din_697), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(o8_status));
SDFFN u15_crac_din_reg_b9_b (.CK(clk_i), .D(n_1028), .Q(crac_din_700), .SO(crac_din_700), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_din_697));
SDFFN u15_crac_din_reg_b12_b (.CK(clk_i), .D(n_1193), .Q(crac_din_703), .SO(crac_din_703), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_din_700));
SDFFN u15_crac_din_reg_b1_b (.CK(clk_i), .D(n_1202), .Q(crac_din_692), .SO(crac_din_692), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_din_703));
SDFFN u15_crac_din_reg_b7_b (.CK(clk_i), .D(n_1022), .Q(crac_din_698), .SO(crac_din_698), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_din_692));
SDFFN u15_crac_din_reg_b14_b (.CK(clk_i), .D(n_1030), .Q(crac_din_705), .SO(crac_din_705), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_din_698));
SDFFN u15_crac_din_reg_b10_b (.CK(clk_i), .D(n_1031), .Q(crac_din_701), .SO(crac_din_701), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_din_705));
SDFFN u15_crac_din_reg_b15_b (.CK(clk_i), .D(n_1083), .Q(crac_din_706), .SO(crac_din_706), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_din_701));
SDFFN u15_crac_din_reg_b4_b (.CK(clk_i), .D(n_1034), .Q(crac_din_695), .SO(crac_din_695), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_din_706));
SDFFN u15_crac_din_reg_b8_b (.CK(clk_i), .D(n_1037), .Q(crac_din_699), .SO(crac_din_699), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_din_695));
SDFFN u15_crac_din_reg_b11_b (.CK(clk_i), .D(n_1029), .Q(crac_din_702), .SO(crac_din_702), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_din_699));
SDFFN u15_crac_din_reg_b13_b (.CK(clk_i), .D(n_1192), .Q(crac_din_704), .SO(crac_din_704), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_din_702));
SDFFN u15_crac_din_reg_b2_b (.CK(clk_i), .D(n_1194), .Q(crac_din_693), .SO(crac_din_693), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_din_704));
SDFFN u15_crac_din_reg_b0_b (.CK(clk_i), .D(n_1074), .Q(crac_din), .SO(crac_din), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_din_693));
SDFFN u15_crac_din_reg_b5_b (.CK(clk_i), .D(n_1197), .Q(crac_din_696), .SO(crac_din_696), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(crac_din));
SDFFNSRN u5_status_reg_b0_b (.CK(clk_i), .D(n_6047), .Q(o6_status), .SO(o6_status), .SE(scan_enable), .SI(crac_din_696));
SDFFNSRN u8_status_reg_b0_b (.CK(clk_i), .D(n_5622), .Q(o9_status), .SO(o9_status), .SE(scan_enable), .SI(o6_status));
SDFFN u15_crac_din_reg_b3_b (.CK(clk_i), .D(n_1047), .Q(crac_din_694), .SO(crac_din_694), .RT(1'b0), .ST(1'b0), .SE(scan_enable), .SI(o9_status));
SDFFNSRN u12_we2_reg (.CK(clk_i), .D(n_870), .Q(u12_we2), .SO(u12_we2), .SE(scan_enable), .SI(crac_din_694));
SDFFNSRN u2_bit_clk_r1_reg (.CK(clk_i), .D(n_719), .Q(u2_bit_clk_r1), .SO(u2_bit_clk_r1), .SE(scan_enable), .SI(u12_we2));
SDFFNSRN u12_dout_reg_b7_b (.CK(clk_i), .D(wb_data_i_b7_b), .Q(wb_din_667), .SO(wb_din_667), .SE(scan_enable), .SI(u2_bit_clk_r1));
SDFFNSRN u12_dout_reg_b4_b (.CK(clk_i), .D(wb_data_i_b4_b), .Q(wb_din_664), .SO(wb_din_664), .SE(scan_enable), .SI(wb_din_667));
SDFFNSRN u12_dout_reg_b12_b (.CK(clk_i), .D(wb_data_i_b12_b), .Q(wb_din_672), .SO(wb_din_672), .SE(scan_enable), .SI(wb_din_664));
SDFFNSRN u12_dout_reg_b24_b (.CK(clk_i), .D(wb_data_i_b24_b), .Q(wb_din_684), .SO(wb_din_684), .SE(scan_enable), .SI(wb_din_672));
SDFFNSRN u12_dout_reg_b26_b (.CK(clk_i), .D(wb_data_i_b26_b), .Q(wb_din_686), .SO(wb_din_686), .SE(scan_enable), .SI(wb_din_684));
SDFFNSRN u12_dout_reg_b23_b (.CK(clk_i), .D(wb_data_i_b23_b), .Q(wb_din_683), .SO(wb_din_683), .SE(scan_enable), .SI(wb_din_686));
SDFFNSRN u12_dout_reg_b11_b (.CK(clk_i), .D(wb_data_i_b11_b), .Q(wb_din_671), .SO(wb_din_671), .SE(scan_enable), .SI(wb_din_683));
SDFFNSRN u12_dout_reg_b31_b (.CK(clk_i), .D(wb_data_i_b31_b), .Q(wb_din_691), .SO(wb_din_691), .SE(scan_enable), .SI(wb_din_671));
SDFFNSRN u12_dout_reg_b13_b (.CK(clk_i), .D(wb_data_i_b13_b), .Q(wb_din_673), .SO(wb_din_673), .SE(scan_enable), .SI(wb_din_691));
SDFFNSRN u12_dout_reg_b29_b (.CK(clk_i), .D(wb_data_i_b29_b), .Q(wb_din_689), .SO(wb_din_689), .SE(scan_enable), .SI(wb_din_673));
SDFFNSRN u12_dout_reg_b22_b (.CK(clk_i), .D(wb_data_i_b22_b), .Q(wb_din_682), .SO(wb_din_682), .SE(scan_enable), .SI(wb_din_689));
SDFFNSRN u12_dout_reg_b30_b (.CK(clk_i), .D(wb_data_i_b30_b), .Q(wb_din_690), .SO(wb_din_690), .SE(scan_enable), .SI(wb_din_682));
SDFFNSRN u12_dout_reg_b15_b (.CK(clk_i), .D(wb_data_i_b15_b), .Q(wb_din_675), .SO(wb_din_675), .SE(scan_enable), .SI(wb_din_690));
SDFFNSRN u12_dout_reg_b19_b (.CK(clk_i), .D(wb_data_i_b19_b), .Q(wb_din_679), .SO(wb_din_679), .SE(scan_enable), .SI(wb_din_675));
SDFFNSRN u2_bit_clk_r_reg (.CK(clk_i), .D(bit_clk_pad_i), .Q(u2_bit_clk_r), .SO(u2_bit_clk_r), .SE(scan_enable), .SI(wb_din_679));
SDFFNSRN u12_dout_reg_b27_b (.CK(clk_i), .D(wb_data_i_b27_b), .Q(wb_din_687), .SO(wb_din_687), .SE(scan_enable), .SI(u2_bit_clk_r));
SDFFNSRN u12_dout_reg_b28_b (.CK(clk_i), .D(wb_data_i_b28_b), .Q(wb_din_688), .SO(wb_din_688), .SE(scan_enable), .SI(wb_din_687));
SDFFNSRN u12_dout_reg_b10_b (.CK(clk_i), .D(wb_data_i_b10_b), .Q(wb_din_670), .SO(wb_din_670), .SE(scan_enable), .SI(wb_din_688));
SDFFNSRN u12_dout_reg_b6_b (.CK(clk_i), .D(wb_data_i_b6_b), .Q(wb_din_666), .SO(wb_din_666), .SE(scan_enable), .SI(wb_din_670));
SDFFNSRN u12_dout_reg_b20_b (.CK(clk_i), .D(wb_data_i_b20_b), .Q(wb_din_680), .SO(wb_din_680), .SE(scan_enable), .SI(wb_din_666));
SDFFNSRN u12_dout_reg_b0_b (.CK(clk_i), .D(wb_data_i_b0_b), .Q(wb_din), .SO(wb_din), .SE(scan_enable), .SI(wb_din_680));
SDFFNSRN u12_dout_reg_b21_b (.CK(clk_i), .D(wb_data_i_b21_b), .Q(wb_din_681), .SO(wb_din_681), .SE(scan_enable), .SI(wb_din));
SDFFNSRN u12_dout_reg_b5_b (.CK(clk_i), .D(wb_data_i_b5_b), .Q(wb_din_665), .SO(wb_din_665), .SE(scan_enable), .SI(wb_din_681));
SDFFNSRN u12_dout_reg_b18_b (.CK(clk_i), .D(wb_data_i_b18_b), .Q(wb_din_678), .SO(wb_din_678), .SE(scan_enable), .SI(wb_din_665));
SDFFNSRN u12_dout_reg_b25_b (.CK(clk_i), .D(wb_data_i_b25_b), .Q(wb_din_685), .SO(wb_din_685), .SE(scan_enable), .SI(wb_din_678));
SDFFNSRN u12_dout_reg_b2_b (.CK(clk_i), .D(wb_data_i_b2_b), .Q(wb_din_662), .SO(wb_din_662), .SE(scan_enable), .SI(wb_din_685));
SDFFNSRN u12_dout_reg_b9_b (.CK(clk_i), .D(wb_data_i_b9_b), .Q(wb_din_669), .SO(wb_din_669), .SE(scan_enable), .SI(wb_din_662));
SDFFNSRN u12_dout_reg_b17_b (.CK(clk_i), .D(wb_data_i_b17_b), .Q(wb_din_677), .SO(wb_din_677), .SE(scan_enable), .SI(wb_din_669));
SDFFNSRN u12_dout_reg_b3_b (.CK(clk_i), .D(wb_data_i_b3_b), .Q(wb_din_663), .SO(wb_din_663), .SE(scan_enable), .SI(wb_din_677));
SDFFNSRN u12_dout_reg_b8_b (.CK(clk_i), .D(wb_data_i_b8_b), .Q(wb_din_668), .SO(wb_din_668), .SE(scan_enable), .SI(wb_din_663));
SDFFNSRN u12_dout_reg_b16_b (.CK(clk_i), .D(wb_data_i_b16_b), .Q(wb_din_676), .SO(wb_din_676), .SE(scan_enable), .SI(wb_din_668));
SDFFNSRN u12_dout_reg_b14_b (.CK(clk_i), .D(wb_data_i_b14_b), .Q(wb_din_674), .SO(wb_din_674), .SE(scan_enable), .SI(wb_din_676));
SDFFNSRN u12_dout_reg_b1_b (.CK(clk_i), .D(wb_data_i_b1_b), .Q(wb_din_661), .SO(wb_din_661), .SE(scan_enable), .SI(wb_din_674));
// scan chain ends here

 buf1 BUFbread(scan_data_out, wb_din_661);
NAND2X1 g34356(.A (u8_mem_b3_b_122 ), .B (n_7976), .Y (n_8047));
NAND2X1 g40697(.A (n_715), .B (u15_rdd3), .Y (n_716));
NAND2X1 g31726(.A (n_5502), .B (n_10376), .Y (n_10349));
NAND2X1 g34357(.A (u4_mem_b1_b_75 ), .B (n_7984), .Y (n_8046));
INVX2 g40546(.A (wb_din_690), .Y (n_2864));
NAND2X1 g37737(.A (n_3264), .B (n_2889), .Y (n_4599));
AOI22X1 g37736(.A0 (n_379), .A1 (n_2544), .B0 (n_5359), .B1 (n_1316),.Y (n_1675));
NAND2X1 g37735(.A (n_2404), .B (n_2250), .Y (n_3917));
AOI22X1 g37734(.A0 (n_2558), .A1 (n_1677), .B0 (n_1676), .B1(n_1839), .Y (n_1678));
AOI22X1 g37733(.A0 (n_2502), .A1 (n_1680), .B0 (n_1679), .B1(n_1859), .Y (n_1681));
AOI22X1 g37732(.A0 (n_147), .A1 (n_940), .B0 (n_5512), .B1 (n_1316),.Y (n_2548));
AOI22X1 g37731(.A0 (n_2558), .A1 (n_2550), .B0 (n_2549), .B1(n_2534), .Y (n_2551));
NAND2X1 g37730(.A (n_1523), .B (n_4234), .Y (n_5215));
NAND2X1 g37739(.A (n_2444), .B (n_2320), .Y (n_3916));
AOI22X1 g37738(.A0 (n_143), .A1 (n_2530), .B0 (n_2627), .B1 (n_2544),.Y (n_2628));
OAI21X1 g33027(.A0 (n_7251), .A1 (n_7188), .B0 (n_10518), .Y(n_11974));
OAI21X1 g33026(.A0 (n_7314), .A1 (n_7094), .B0 (n_10518), .Y(n_11990));
OAI21X1 g33025(.A0 (n_7253), .A1 (n_7016), .B0 (n_10518), .Y(n_11954));
OAI21X1 g33024(.A0 (n_7315), .A1 (n_7189), .B0 (n_10518), .Y(n_11978));
OAI21X1 g33023(.A0 (n_7316), .A1 (n_6918), .B0 (n_10518), .Y(n_11952));
OAI21X1 g33022(.A0 (n_7254), .A1 (n_7190), .B0 (n_10518), .Y(n_11968));
OAI21X1 g33021(.A0 (n_7255), .A1 (n_7192), .B0 (n_10518), .Y(n_11970));
OAI21X1 g33020(.A0 (n_7257), .A1 (n_7193), .B0 (n_10518), .Y(n_11964));
MX2X1 g37221(.A (u9_mem_b1_b_143 ), .B (n_4755), .S0 (n_4783), .Y(n_4788));
MX2X1 g37220(.A (u9_mem_b1_b_141 ), .B (n_4757), .S0 (n_4783), .Y(n_4789));
MX2X1 g37223(.A (u9_mem_b1_b_146 ), .B (n_4772), .S0 (n_4783), .Y(n_4785));
MX2X1 g37225(.A (u9_mem_b1_b_148 ), .B (n_4764), .S0 (n_4783), .Y(n_4782));
MX2X1 g37224(.A (u9_mem_b1_b_147 ), .B (n_4769), .S0 (n_4783), .Y(n_4784));
OAI21X1 g33029(.A0 (n_7249), .A1 (n_7186), .B0 (n_10518), .Y(n_11972));
OAI21X1 g33028(.A0 (n_7250), .A1 (n_7093), .B0 (n_10518), .Y(n_10523));
INVX1 g42641(.A (n_1819), .Y (n_742));
MX2X1 g33140(.A (wb_din_672), .B (n_8567), .S0 (n_8538), .Y (n_8568));
NAND2X1 g34353(.A (u4_mem_b1_b_72 ), .B (n_7984), .Y (n_8051));
MX2X1 g33145(.A (wb_din_677), .B (oc2_cfg_984), .S0 (n_8538), .Y(n_8560));
AOI21X1 g40384(.A0 (u26_ps_cnt_b1_b ), .A1 (n_529), .B0 (n_819), .Y(n_1441));
AND2X1 g41518(.A (n_627), .B (n_626), .Y (n_858));
XOR2X1 g40385(.A (u8_wp_b1_b ), .B (n_12280), .Y (n_1929));
MX2X1 g36176(.A (n_6349), .B (n_6486), .S0 (n_6359), .Y (n_6350));
MX2X1 g36177(.A (n_6347), .B (n_6547), .S0 (n_6359), .Y (n_6348));
MX2X1 g36174(.A (n_6353), .B (n_6442), .S0 (n_6359), .Y (n_6354));
MX2X1 g36175(.A (n_6351), .B (n_6544), .S0 (n_6359), .Y (n_6352));
MX2X1 g36172(.A (n_6357), .B (n_6497), .S0 (n_6359), .Y (n_6358));
MX2X1 g36173(.A (n_6355), .B (n_6444), .S0 (n_6359), .Y (n_6356));
MX2X1 g36171(.A (n_5949), .B (n_6008), .S0 (n_6341), .Y (n_5950));
NAND2X1 g38853(.A (u5_mem_b3_b_136 ), .B (n_1543), .Y (n_1333));
MX2X1 g36178(.A (n_6344), .B (n_6483), .S0 (n_6359), .Y (n_6345));
MX2X1 g36179(.A (n_5947), .B (n_5983), .S0 (n_6359), .Y (n_5948));
INVX1 g42702(.A (u10_mem_b2_b_108 ), .Y (n_39));
NAND2X1 g39025(.A (n_12826), .B (u3_mem_b0_b_108 ), .Y (n_3502));
INVX1 g42700(.A (u9_mem_b1_b_124 ), .Y (n_6942));
INVX1 g42706(.A (n_862), .Y (n_11043));
AOI22X1 g40382(.A0 (n_494), .A1 (n_1446), .B0 (u8_rp_b3_b ), .B1(u8_wp_b2_b ), .Y (n_1447));
AOI21X1 g35565(.A0 (n_6818), .A1 (n_6135), .B0 (n_12145), .Y(n_7328));
AOI21X1 g35566(.A0 (n_6313), .A1 (n_6133), .B0 (n_7324), .Y (n_7278));
INVX1 g31771(.A (n_9604), .Y (n_9605));
AOI21X1 g31770(.A0 (n_1208), .A1 (n_7160), .B0 (n_9503), .Y (n_9554));
INVX1 g31773(.A (n_9552), .Y (n_9553));
AOI21X1 g31772(.A0 (n_1071), .A1 (n_7036), .B0 (n_9560), .Y (n_9604));
INVX1 g31775(.A (n_9550), .Y (n_9551));
AOI21X1 g31774(.A0 (n_1130), .A1 (n_7035), .B0 (n_9501), .Y (n_9552));
AOI21X1 g31777(.A0 (n_8847), .A1 (n_7532), .B0 (n_7527), .Y (n_8848));
AOI21X1 g31776(.A0 (n_1116), .A1 (n_7034), .B0 (n_9499), .Y (n_9550));
AOI21X1 g31779(.A0 (n_9444), .A1 (n_8208), .B0 (n_8206), .Y (n_9445));
AOI21X1 g31778(.A0 (n_8843), .A1 (n_7529), .B0 (n_7525), .Y (n_8844));
INVX4 g45473(.A (n_12357), .Y (n_11934));
NAND2X1 g39020(.A (u6_mem_b2_b_45 ), .B (n_3474), .Y (n_3509));
AOI21X1 g35850(.A0 (n_2583), .A1 (n_4716), .B0 (n_7353), .Y (n_7108));
NOR2X1 g35851(.A (n_4665), .B (n_7353), .Y (n_7107));
NOR2X1 g35852(.A (n_4662), .B (n_7353), .Y (n_7151));
NOR2X1 g35853(.A (n_1292), .B (n_4104), .Y (n_4105));
AOI21X1 g35678(.A0 (n_877), .A1 (n_1221), .B0 (i3_re), .Y (n_6708));
AOI21X1 g35679(.A0 (n_1232), .A1 (n_2364), .B0 (i4_re), .Y (n_6707));
AOI21X1 g30828(.A0 (n_11964), .A1 (n_11965), .B0 (n_11086), .Y(n_11095));
AOI21X1 g30829(.A0 (n_11970), .A1 (n_11971), .B0 (n_5827), .Y(n_11094));
AOI21X1 g30826(.A0 (n_9915), .A1 (n_9798), .B0 (n_10916), .Y(n_10909));
AOI21X1 g30827(.A0 (n_9914), .A1 (n_9797), .B0 (n_2485), .Y(n_10908));
AOI21X1 g30824(.A0 (n_12813), .A1 (n_12814), .B0 (n_2485), .Y(n_10911));
AOI21X1 g30825(.A0 (n_12815), .A1 (n_12816), .B0 (n_10916), .Y(n_10910));
AOI21X1 g30822(.A0 (n_12610), .A1 (n_11999), .B0 (n_10921), .Y(n_10913));
AOI21X1 g30823(.A0 (n_12811), .A1 (n_12812), .B0 (n_2485), .Y(n_10912));
NOR2X1 g30820(.A (n_10786), .B (n_10994), .Y (n_10996));
NOR2X1 g30821(.A (n_10784), .B (n_10994), .Y (n_10995));
INVX2 g45689(.A (n_12384), .Y (n_12385));
CLKBUFX1 g41732(.A (n_1040), .Y (n_2513));
INVX4 g45692(.A (n_12385), .Y (n_12389));
NAND2X1 g39432(.A (n_1068), .B (u7_rp_b3_b ), .Y (n_4080));
INVX1 g37001(.A (n_6226), .Y (n_5702));
MX2X1 g38760(.A (u3_mem_b0_b_94 ), .B (wb_din_664), .S0 (n_3807), .Y(n_3575));
NAND2X1 g39479(.A (u6_mem_b1_b_64 ), .B (n_4253), .Y (n_11712));
MX2X1 g38763(.A (u3_mem_b0_b_98 ), .B (wb_din_668), .S0 (n_3807), .Y(n_3572));
NOR2X1 g35569(.A (n_1080), .B (i6_re), .Y (n_6715));
NAND2X1 g39476(.A (n_11798), .B (u8_mem_b0_b_105 ), .Y (n_11461));
MX2X1 g38762(.A (u6_mem_b0_b_109 ), .B (wb_din_679), .S0 (n_3632), .Y(n_3573));
AOI21X1 g35553(.A0 (n_5592), .A1 (n_4731), .B0 (n_7353), .Y (n_7140));
NAND2X1 g39433(.A (u4_mem_b1_b_61 ), .B (n_12259), .Y (n_4192));
NAND2X1 g39474(.A (u6_mem_b1_b_65 ), .B (n_12169), .Y (n_11714));
MX2X1 g38764(.A (u7_mem_b0_b_115 ), .B (wb_din_685), .S0 (n_3622), .Y(n_3571));
NAND2X1 g39779(.A (u7_mem_b2_b_52 ), .B (n_12650), .Y (n_4128));
NOR2X1 g39778(.A (n_3332), .B (n_2801), .Y (n_2964));
NAND2X1 g39770(.A (u7_mem_b2_b_35 ), .B (n_12654), .Y (n_2969));
NAND2X1 g39773(.A (n_2302), .B (in_slt_434), .Y (n_4751));
MX2X1 g38766(.A (u7_mem_b0_b_113 ), .B (wb_din_683), .S0 (n_3622), .Y(n_3569));
NAND2X1 g39775(.A (n_2325), .B (in_slt_447), .Y (n_2249));
NAND2X1 g39774(.A (u7_mem_b2_b_51 ), .B (n_12645), .Y (n_4129));
NOR2X1 g39777(.A (n_4996), .B (n_2720), .Y (n_2965));
NAND2X1 g39776(.A (u7_mem_b2_b_37 ), .B (n_12654), .Y (n_2966));
MX2X1 g38768(.A (u6_mem_b0_b_104 ), .B (wb_din_674), .S0 (n_3632), .Y(n_3567));
NAND2X1 g39430(.A (u7_mem_b2_b_38 ), .B (n_12641), .Y (n_3188));
INVX4 g41739(.A (n_1360), .Y (n_4560));
MX2X1 g31195(.A (n_6481), .B (n_419), .S0 (n_10513), .Y (n_10542));
MX2X1 g31194(.A (n_5985), .B (n_5984), .S0 (n_10513), .Y (n_10543));
MX2X1 g31197(.A (n_6477), .B (n_6476), .S0 (n_10315), .Y (n_10215));
MX2X1 g31196(.A (n_6480), .B (n_6479), .S0 (n_10537), .Y (n_10540));
MX2X1 g31191(.A (n_6549), .B (n_6548), .S0 (n_10537), .Y (n_10546));
MX2X1 g31190(.A (n_6488), .B (n_6487), .S0 (n_10513), .Y (n_10547));
MX2X1 g31193(.A (n_5982), .B (n_5981), .S0 (n_10565), .Y (n_10544));
MX2X1 g31192(.A (n_6485), .B (n_6484), .S0 (n_10537), .Y (n_10545));
MX2X1 g31199(.A (n_6469), .B (n_6468), .S0 (n_10315), .Y (n_10214));
MX2X1 g31198(.A (n_6474), .B (n_433), .S0 (n_10537), .Y (n_10539));
NAND2X1 g38852(.A (u6_mem_b3_b_147 ), .B (n_2465), .Y (n_2440));
OAI21X1 g36701(.A0 (n_5190), .A1 (n_5189), .B0 (n_634), .Y (n_5751));
MX2X1 g34109(.A (u7_mem_b0_b_93 ), .B (n_3616), .S0 (n_7493), .Y(n_8730));
MX2X1 g34108(.A (u7_mem_b0_b_121 ), .B (n_3635), .S0 (n_7493), .Y(n_9393));
MX2X1 g34105(.A (u7_mem_b0_b_119 ), .B (n_3610), .S0 (n_7493), .Y(n_8733));
MX2X1 g34104(.A (u7_mem_b0_b_118 ), .B (n_3636), .S0 (n_7493), .Y(n_8735));
MX2X1 g34107(.A (u7_mem_b0_b_120 ), .B (n_3613), .S0 (n_7493), .Y(n_8731));
MX2X1 g34106(.A (u7_mem_b0_b_92 ), .B (n_3612), .S0 (n_7493), .Y(n_8732));
MX2X1 g34101(.A (u7_mem_b0_b_115 ), .B (n_3571), .S0 (n_7493), .Y(n_8738));
MX2X1 g34100(.A (u7_mem_b0_b_114 ), .B (n_3639), .S0 (n_7493), .Y(n_9394));
MX2X1 g34103(.A (u7_mem_b0_b_117 ), .B (n_3607), .S0 (n_7493), .Y(n_8736));
MX2X1 g34102(.A (u7_mem_b0_b_116 ), .B (n_3638), .S0 (n_7493), .Y(n_8737));
AOI21X1 g35557(.A0 (n_5589), .A1 (n_4724), .B0 (n_7353), .Y (n_7136));
NAND2X1 g39087(.A (n_4560), .B (in_slt_450), .Y (n_5315));
NAND2X1 g36356(.A (n_6821), .B (n_5844), .Y (n_5920));
NAND2X1 g39085(.A (n_11804), .B (u8_mem_b0_b_113 ), .Y (n_3460));
NAND2X1 g39084(.A (u5_mem_b2_b_42 ), .B (n_12823), .Y (n_12806));
NOR2X1 g39083(.A (n_2691), .B (n_1488), .Y (n_1501));
NOR2X1 g39082(.A (n_3089), .B (n_3008), .Y (n_3463));
NOR2X1 g39081(.A (n_5138), .B (n_2702), .Y (n_3465));
NAND2X1 g39080(.A (in_slt_413), .B (n_3415), .Y (n_3466));
OR2X1 g36354(.A (n_2617), .B (n_3944), .Y (n_2618));
NAND2X1 g39088(.A (n_11798), .B (u8_mem_b0_b_100 ), .Y (n_11451));
OAI21X1 g33597(.A0 (n_5072), .A1 (n_9349), .B0 (n_7955), .Y (n_9325));
OAI21X1 g33596(.A0 (n_5074), .A1 (n_9326), .B0 (n_7956), .Y (n_9327));
OAI21X1 g33595(.A0 (n_5075), .A1 (n_9326), .B0 (n_7958), .Y (n_9328));
OAI21X1 g33594(.A0 (n_5077), .A1 (n_9336), .B0 (n_7959), .Y (n_9329));
OAI21X1 g33592(.A0 (n_5080), .A1 (n_9333), .B0 (n_7961), .Y (n_9331));
OAI21X1 g33591(.A0 (n_5081), .A1 (n_9333), .B0 (n_7962), .Y (n_9332));
OAI21X1 g33590(.A0 (n_5082), .A1 (n_9333), .B0 (n_7963), .Y (n_9334));
NOR2X1 g40246(.A (n_2780), .B (n_2729), .Y (n_2695));
NAND2X1 g36352(.A (n_6821), .B (n_5851), .Y (n_5922));
OAI21X1 g33599(.A0 (n_5068), .A1 (n_9326), .B0 (n_7953), .Y (n_9322));
OAI21X1 g33598(.A0 (n_5071), .A1 (n_9349), .B0 (n_7954), .Y (n_9324));
OAI21X1 g33849(.A0 (n_4466), .A1 (n_9055), .B0 (n_7675), .Y (n_9009));
OAI21X1 g33848(.A0 (n_4314), .A1 (n_9010), .B0 (n_7676), .Y (n_9011));
NAND2X1 g36350(.A (n_5853), .B (n_6821), .Y (n_5923));
OAI21X1 g33841(.A0 (n_4406), .A1 (n_9043), .B0 (n_7683), .Y (n_9019));
OAI21X1 g33840(.A0 (n_4404), .A1 (n_9034), .B0 (n_7684), .Y (n_9020));
OAI21X1 g33843(.A0 (n_4424), .A1 (n_9055), .B0 (n_7681), .Y (n_9016));
OAI21X1 g33842(.A0 (n_4318), .A1 (n_9055), .B0 (n_7682), .Y (n_9018));
OAI21X1 g33845(.A0 (n_4316), .A1 (n_9055), .B0 (n_7679), .Y (n_9014));
OAI21X1 g33844(.A0 (n_4317), .A1 (n_9043), .B0 (n_7680), .Y (n_9015));
OAI21X1 g33847(.A0 (n_4452), .A1 (n_9055), .B0 (n_7677), .Y (n_9012));
OAI21X1 g33846(.A0 (n_4315), .A1 (n_9038), .B0 (n_7678), .Y (n_9013));
MX2X1 g37229(.A (u9_mem_b2_b_109 ), .B (n_4776), .S0 (n_5732), .Y(n_4777));
INVX2 g34968(.A (n_7428), .Y (n_9161));
MX2X1 g37228(.A (u9_mem_b2_b_107 ), .B (n_4778), .S0 (n_6898), .Y(n_4779));
NOR2X1 g39435(.A (n_2712), .B (n_1488), .Y (n_1480));
AOI22X1 g37779(.A0 (n_1756), .A1 (n_6360), .B0 (n_6503), .B1(n_1643), .Y (n_1660));
OR2X1 g38901(.A (n_393), .B (n_2513), .Y (n_2412));
NAND2X1 g38903(.A (u8_mem_b3_b_149 ), .B (n_2468), .Y (n_2410));
MX2X1 g37222(.A (u9_mem_b1_b_145 ), .B (n_4743), .S0 (n_4783), .Y(n_4786));
NAND2X1 g38905(.A (u5_mem_b3_b_122 ), .B (n_3543), .Y (n_2408));
NAND2X1 g38904(.A (u3_mem_b3_b_141 ), .B (n_2463), .Y (n_2409));
MX2X1 g37227(.A (u10_mem_b1_b_145 ), .B (n_4759), .S0 (n_5407), .Y(n_4780));
MX2X1 g37226(.A (u9_mem_b1_b_149 ), .B (n_4767), .S0 (n_5730), .Y(n_4781));
OR2X1 g32645(.A (u11_wp_b0_b ), .B (n_9631), .Y (n_9750));
NAND2X1 g32646(.A (n_9931), .B (n_9833), .Y (n_10949));
NAND2X1 g32647(.A (n_290), .B (n_9931), .Y (n_9933));
NAND2X1 g32640(.A (u10_wp_b3_b ), .B (n_9564), .Y (n_9751));
INVX1 g45441(.A (n_11827), .Y (n_11823));
NAND3X1 g45910(.A (n_12636), .B (n_12634), .C (n_5818), .Y (n_12638));
INVX4 g32643(.A (n_9750), .Y (n_10103));
NAND2X1 g32648(.A (n_287), .B (n_9931), .Y (n_9932));
NAND2X1 g32649(.A (n_84), .B (n_9931), .Y (n_9930));
INVX4 g45919(.A (n_12659), .Y (n_12654));
AOI21X1 g40393(.A0 (u11_rp_b0_b ), .A1 (u11_wp_b1_b ), .B0 (n_916), .Y(n_5442));
XOR2X1 g40391(.A (n_1198), .B (u8_wp_b0_b ), .Y (n_5622));
AOI21X1 g40390(.A0 (n_1206), .A1 (n_5420), .B0 (n_1207), .Y (n_4104));
XOR2X1 g40397(.A (n_1419), .B (n_1923), .Y (n_6049));
AOI21X1 g40396(.A0 (u10_rp_b2_b ), .A1 (u10_wp_b3_b ), .B0 (n_514), .Y(n_1290));
XOR2X1 g40395(.A (n_1421), .B (n_1921), .Y (n_5616));
AOI21X1 g40394(.A0 (u3_rp_b3_b ), .A1 (u3_wp_b2_b ), .B0 (n_477), .Y(n_822));
XOR2X1 g40399(.A (n_6841), .B (n_907), .Y (n_1926));
AOI21X1 g40398(.A0 (u11_rp_b2_b ), .A1 (u11_wp_b3_b ), .B0 (n_522), .Y(n_2617));
MX2X1 g38758(.A (u3_mem_b0_b_121 ), .B (wb_din_691), .S0 (n_3807), .Y(n_3577));
MX2X1 g38759(.A (u6_mem_b0_b_107 ), .B (wb_din_677), .S0 (n_3632), .Y(n_3576));
XOR2X1 g38028(.A (u11_wp_b3_b ), .B (n_695), .Y (n_1025));
AOI21X1 g38029(.A0 (u3_mem_b1_b_72 ), .A1 (n_5148), .B0 (n_2677), .Y(n_5143));
NAND4X1 g37034(.A (n_4127), .B (n_2294), .C (n_3120), .D (n_1530), .Y(n_6211));
INVX1 g37035(.A (n_6233), .Y (n_5690));
NAND4X1 g37036(.A (n_4173), .B (n_2959), .C (n_3093), .D (n_1537), .Y(n_6233));
NAND4X1 g37037(.A (n_3489), .B (n_3502), .C (n_2898), .D (n_2405), .Y(n_6186));
INVX1 g37030(.A (n_5544), .Y (n_5545));
AOI21X1 g38023(.A0 (u8_mem_b3_b ), .A1 (n_3879), .B0 (n_1503), .Y(n_3886));
NAND4X1 g37032(.A (n_2966), .B (n_3105), .C (n_2493), .D (n_1526), .Y(n_5544));
INVX1 g37033(.A (n_6211), .Y (n_5691));
INVX1 g42359(.A (u10_mem_b0_b_154 ), .Y (n_6335));
OAI21X1 g36619(.A0 (n_4576), .A1 (n_5203), .B0 (n_784), .Y (n_6138));
NAND2X1 g36618(.A (n_5252), .B (n_3980), .Y (n_5795));
NAND2X1 g36349(.A (n_6779), .B (n_6821), .Y (n_6823));
NAND2X1 g36348(.A (n_5855), .B (n_6821), .Y (n_5924));
NAND2X1 g36345(.A (n_5833), .B (n_6821), .Y (n_5925));
NAND2X1 g36344(.A (n_5835), .B (n_6821), .Y (n_5926));
NAND2X1 g36347(.A (n_12746), .B (n_6824), .Y (n_6825));
NAND2X1 g36346(.A (n_6237), .B (n_6824), .Y (n_6309));
NAND3X1 g36617(.A (n_1284), .B (u12_we2), .C (u12_we1), .Y (n_5248));
NAND2X1 g36340(.A (n_6252), .B (n_6824), .Y (n_6312));
OAI21X1 g36615(.A0 (n_5185), .A1 (n_5184), .B0 (n_634), .Y (n_5796));
NAND2X1 g45708(.A (n_1546), .B (u7_mem_b3_b_140 ), .Y (n_12405));
INVX2 g45591(.A (n_12384), .Y (n_12244));
INVX1 g45703(.A (u5_rp_b1_b ), .Y (n_12400));
INVX1 g45702(.A (n_12581), .Y (n_12399));
NAND2X2 g45701(.A (n_12399), .B (n_12400), .Y (n_12401));
NAND2X1 g45707(.A (n_2491), .B (u7_mem_b0_b_109 ), .Y (n_12404));
NAND2X1 g45706(.A (n_4225), .B (u7_mem_b1_b_78 ), .Y (n_12403));
NAND4X1 g45705(.A (n_12403), .B (n_12404), .C (n_12405), .D(n_12410), .Y (n_12411));
CLKBUFX1 g45704(.A (n_12400), .Y (n_1033));
NOR2X1 g39612(.A (n_3117), .B (n_2686), .Y (n_3058));
INVX2 g40486(.A (wb_din_689), .Y (n_3008));
NAND2X1 g38950(.A (u7_mem_b3_b_141 ), .B (n_1546), .Y (n_1516));
AOI22X1 g37690(.A0 (n_6942), .A1 (n_1859), .B0 (n_6900), .B1(n_1835), .Y (n_1694));
AOI22X1 g37692(.A0 (n_2502), .A1 (n_6849), .B0 (n_6886), .B1(n_1760), .Y (n_1693));
NAND2X1 g37693(.A (n_3531), .B (n_3367), .Y (n_4607));
NAND2X1 g37694(.A (n_4140), .B (n_3366), .Y (n_5219));
AOI22X1 g37695(.A0 (n_6033), .A1 (n_2544), .B0 (n_6013), .B1(n_1316), .Y (n_1692));
NAND2X1 g37697(.A (n_4219), .B (n_3362), .Y (n_5218));
AOI21X1 g37698(.A0 (n_6030), .A1 (n_2553), .B0 (n_2365), .Y (n_4078));
AOI22X1 g37699(.A0 (n_2558), .A1 (n_5955), .B0 (n_6010), .B1(n_1316), .Y (n_1249));
INVX2 g45594(.A (n_12258), .Y (n_12252));
NOR2X1 g41374(.A (n_685), .B (n_708), .Y (n_686));
NOR2X1 g41372(.A (n_8550), .B (oc2_cfg_987), .Y (n_9611));
NOR2X1 g41370(.A (u10_wp_b1_b ), .B (u10_wp_b2_b ), .Y (n_1064));
NOR2X1 g41371(.A (u13_ints_r_b27_b ), .B (ic2_int_set_723), .Y(n_513));
INVX4 g45905(.A (u7_rp_b0_b ), .Y (n_12634));
MX2X1 g31348(.A (u10_din_tmp_44), .B (in_slt_425), .S0 (n_9860), .Y(n_9871));
MX2X1 g31349(.A (u10_din_tmp_45), .B (in_slt_426), .S0 (n_9860), .Y(n_9869));
NAND2X1 g31698(.A (n_298), .B (n_10376), .Y (n_10364));
NAND2X1 g31699(.A (n_236), .B (n_10376), .Y (n_10363));
NOR2X1 g40312(.A (n_2144), .B (n_2755), .Y (n_1968));
NAND2X1 g31692(.A (n_279), .B (n_10376), .Y (n_10369));
NOR2X1 g31693(.A (n_11890), .B (n_1184), .Y (n_9989));
NAND2X1 g31690(.A (n_81), .B (n_10385), .Y (n_10371));
NAND2X1 g31691(.A (n_1627), .B (n_10376), .Y (n_10370));
NAND2X1 g31696(.A (n_270), .B (n_10385), .Y (n_10365));
MX2X1 g31345(.A (n_5963), .B (n_5962), .S0 (n_10137), .Y (n_10118));
XOR2X1 g31346(.A (u7_rp_b0_b ), .B (n_9901), .Y (n_10810));
NAND2X1 g31695(.A (n_275), .B (n_10376), .Y (n_10366));
NAND2X1 g37968(.A (n_2867), .B (n_2876), .Y (n_5175));
NAND2X1 g37969(.A (n_1812), .B (n_3442), .Y (n_5174));
AOI22X1 g37962(.A0 (n_6457), .A1 (n_940), .B0 (n_6591), .B1 (n_1316),.Y (n_3892));
NAND2X1 g37963(.A (n_3419), .B (n_3460), .Y (n_5178));
NAND2X1 g37960(.A (n_3003), .B (n_3429), .Y (n_5180));
NAND2X1 g37961(.A (n_2396), .B (n_2844), .Y (n_5179));
NAND2X1 g37966(.A (n_2852), .B (n_3160), .Y (n_5176));
NAND2X1 g37967(.A (n_2383), .B (n_2301), .Y (n_4552));
NAND2X1 g37964(.A (n_2375), .B (n_2891), .Y (n_5177));
AOI22X1 g37965(.A0 (n_2502), .A1 (n_6394), .B0 (n_6537), .B1(n_1859), .Y (n_2503));
NAND2X1 g33278(.A (u15_rdd1), .B (n_9688), .Y (n_9795));
NAND2X1 g33279(.A (crac_wr), .B (n_9689), .Y (n_9794));
INVX1 g33272(.A (n_9571), .Y (n_9631));
NOR2X1 g33273(.A (n_8210), .B (u14_u8_en_out_l2), .Y (n_9571));
NAND2X1 g39339(.A (u5_mem_b1_b_81 ), .B (n_3239), .Y (n_3264));
NOR2X1 g33277(.A (n_9711), .B (n_294), .Y (n_9712));
NAND3X1 g33274(.A (n_991), .B (n_614), .C (n_7984), .Y (n_8179));
AND2X1 g33275(.A (n_7521), .B (wb_din_661), .Y (n_7522));
INVX1 g42139(.A (u11_mem_b2_b_95 ), .Y (n_6431));
NOR2X1 g39492(.A (n_2720), .B (n_1488), .Y (n_1272));
NAND3X1 g45907(.A (n_12635), .B (n_12636), .C (u7_rp_b0_b ), .Y(n_12637));
INVX1 g42130(.A (u10_mem_b3_b ), .Y (n_6005));
INVX1 g42137(.A (u9_mem_b0_b_153 ), .Y (n_6854));
NAND2X1 g39338(.A (u6_mem_b2_b_40 ), .B (n_3474), .Y (n_11698));
MX2X1 g35991(.A (n_6483), .B (n_6650), .S0 (n_6649), .Y (n_6651));
MX2X1 g35990(.A (n_6652), .B (n_6579), .S0 (n_5341), .Y (n_6653));
MX2X1 g35993(.A (n_6942), .B (n_6899), .S0 (n_5730), .Y (n_6943));
MX2X1 g35992(.A (n_6945), .B (n_6913), .S0 (n_5730), .Y (n_6946));
MX2X1 g35995(.A (n_6937), .B (n_6906), .S0 (n_4783), .Y (n_6938));
MX2X1 g35994(.A (n_6940), .B (n_6927), .S0 (n_4783), .Y (n_6941));
MX2X1 g35997(.A (n_6644), .B (n_6618), .S0 (n_6898), .Y (n_6645));
MX2X1 g35999(.A (n_6638), .B (n_6637), .S0 (n_6898), .Y (n_6639));
MX2X1 g35998(.A (n_6641), .B (n_6533), .S0 (n_6898), .Y (n_6642));
NOR2X1 g39966(.A (n_704), .B (u2_to_cnt_b1_b ), .Y (n_1051));
NAND2X1 g39967(.A (n_11804), .B (u8_mem_b0_b_91 ), .Y (n_11742));
NAND2X1 g39960(.A (n_11804), .B (u8_mem_b0_b_108 ), .Y (n_3890));
NAND2X1 g39961(.A (n_2325), .B (in_slt_453), .Y (n_2227));
NOR2X1 g39962(.A (n_3089), .B (n_2741), .Y (n_2851));
NAND2X1 g39963(.A (u8_mem_b1_b_77 ), .B (n_12291), .Y (n_2850));
INVX4 g45497(.A (n_12076), .Y (n_12087));
INVX4 g45496(.A (n_12076), .Y (n_12079));
INVX1 g35199(.A (n_7396), .Y (n_8930));
INVX1 g35190(.A (n_7396), .Y (n_8433));
INVX1 g35193(.A (n_7396), .Y (n_8449));
INVX1 g35192(.A (n_7396), .Y (n_8453));
INVX1 g35195(.A (n_7396), .Y (n_8457));
INVX1 g35197(.A (n_7396), .Y (n_8464));
INVX1 g35196(.A (n_7396), .Y (n_8438));
NAND2X1 g34822(.A (u8_mem_b1_b_73 ), .B (n_7976), .Y (n_7612));
NAND2X1 g34823(.A (u8_mem_b1_b_74 ), .B (n_7976), .Y (n_7611));
NAND2X1 g34820(.A (u8_mem_b1_b_70 ), .B (n_7976), .Y (n_7614));
NAND2X1 g34821(.A (u8_mem_b1_b_72 ), .B (n_7976), .Y (n_7613));
NAND2X1 g34826(.A (u8_mem_b1_b_77 ), .B (n_7976), .Y (n_7608));
NAND2X1 g34827(.A (u3_mem_b1_b_90 ), .B (n_8101), .Y (n_7607));
NAND2X1 g34824(.A (u8_mem_b1_b_76 ), .B (n_7976), .Y (n_7610));
NAND2X1 g34825(.A (u8_mem_b3_b_133 ), .B (n_7976), .Y (n_7609));
NAND2X1 g34828(.A (u8_mem_b1_b_78 ), .B (n_7976), .Y (n_7606));
NAND2X1 g34829(.A (u8_mem_b1_b_79 ), .B (n_7976), .Y (n_7605));
NAND3X1 g45903(.A (n_12634), .B (n_12636), .C (n_11855), .Y(n_12631));
AOI21X1 g30123(.A0 (n_6839), .A1 (n_11136), .B0 (n_10960), .Y(n_11142));
AOI21X1 g30122(.A0 (n_6836), .A1 (n_12589), .B0 (n_10963), .Y(n_11526));
AOI22X1 g30121(.A0 (n_9581), .A1 (n_9650), .B0 (n_599), .B1 (n_9499),.Y (n_9753));
AOI22X1 g30120(.A0 (n_9582), .A1 (n_9653), .B0 (n_690), .B1 (n_9501),.Y (n_9754));
AOI21X1 g30127(.A0 (n_6059), .A1 (n_11136), .B0 (n_10959), .Y(n_11505));
NAND2X1 g35446(.A (n_7301), .B (n_6696), .Y (n_7455));
AOI21X1 g30125(.A0 (n_6842), .A1 (n_11126), .B0 (n_11005), .Y(n_11522));
AOI21X1 g30124(.A0 (n_7049), .A1 (n_11131), .B0 (n_11007), .Y(n_11520));
NAND2X1 g39348(.A (n_3255), .B (u5_mem_b0_b_97 ), .Y (n_3256));
NAND2X1 g39349(.A (n_2330), .B (u7_mem_b0_b_91 ), .Y (n_2321));
MX2X1 g30129(.A (n_6756), .B (n_10328), .S0 (n_10985), .Y (n_10970));
MX2X1 g30128(.A (n_7010), .B (n_10330), .S0 (n_10992), .Y (n_10971));
AOI21X1 g35339(.A0 (i4_dout), .A1 (n_7468), .B0 (n_7352), .Y(n_7475));
NOR2X1 g35338(.A (n_5445), .B (u2_bit_clk_e), .Y (n_6054));
NAND4X1 g36978(.A (n_3161), .B (n_2247), .C (n_3514), .D (n_1521), .Y(n_6147));
NAND2X1 g36977(.A (n_1574), .B (n_1573), .Y (n_4004));
INVX1 g36975(.A (n_5833), .Y (n_5553));
NAND4X1 g36972(.A (n_11717), .B (n_11718), .C (n_2286), .D (n_2428),.Y (n_5855));
INVX1 g36973(.A (n_12171), .Y (n_6076));
NAND2X1 g36970(.A (n_1577), .B (n_1576), .Y (n_4005));
INVX1 g36971(.A (n_5855), .Y (n_5554));
CLKBUFX3 g32872(.A (n_9724), .Y (n_10081));
BUFX3 g32871(.A (n_9632), .Y (n_9676));
INVX2 g32875(.A (n_9829), .Y (n_10565));
NAND2X1 g39331(.A (u4_mem_b1_b_82 ), .B (n_12267), .Y (n_4200));
NOR2X1 g40054(.A (n_2169), .B (n_2681), .Y (n_2170));
NOR2X1 g40055(.A (n_2038), .B (n_2786), .Y (n_2168));
NAND2X1 g34311(.A (u3_mem_b3_b_147 ), .B (n_8141), .Y (n_8085));
OAI21X1 g33472(.A0 (n_4871), .A1 (n_9022), .B0 (n_8100), .Y (n_8386));
OAI21X1 g33473(.A0 (n_4889), .A1 (n_8383), .B0 (n_8099), .Y (n_8385));
OAI21X1 g33474(.A0 (n_5139), .A1 (n_8383), .B0 (n_8098), .Y (n_8384));
NAND2X1 g34316(.A (n_6675), .B (n_7459), .Y (n_8244));
OAI21X1 g33477(.A0 (n_5136), .A1 (n_8380), .B0 (n_8094), .Y (n_8379));
OAI21X1 g33478(.A0 (n_5135), .A1 (n_8380), .B0 (n_8093), .Y (n_8378));
OAI21X1 g33479(.A0 (n_4910), .A1 (n_8375), .B0 (n_8092), .Y (n_8377));
INVX1 g37087(.A (n_5898), .Y (n_5534));
NAND2X1 g34648(.A (u6_mem_b2_b_51 ), .B (n_7758), .Y (n_7777));
OAI21X1 g33969(.A0 (n_4434), .A1 (n_8449), .B0 (n_7977), .Y (n_8855));
NAND2X1 g34646(.A (u6_mem_b2_b_49 ), .B (n_7758), .Y (n_7779));
NAND2X1 g34647(.A (u6_mem_b2_b_50 ), .B (n_7758), .Y (n_7778));
NAND2X1 g39335(.A (n_3255), .B (u5_mem_b0_b_96 ), .Y (n_3268));
NAND2X1 g34645(.A (u6_mem_b2_b_48 ), .B (n_7758), .Y (n_7780));
OAI21X1 g33963(.A0 (n_4304), .A1 (n_8891), .B0 (n_7662), .Y (n_8862));
OAI21X1 g33960(.A0 (n_4860), .A1 (n_8856), .B0 (n_7570), .Y (n_8866));
OAI21X1 g33961(.A0 (n_4298), .A1 (n_8868), .B0 (n_7700), .Y (n_8865));
AOI21X1 g38255(.A0 (u6_mem_b3_b_145 ), .A1 (n_5059), .B0 (n_3175), .Y(n_5055));
NAND2X1 g37750(.A (n_3130), .B (n_3231), .Y (n_4594));
XOR2X1 g37201(.A (n_1417), .B (n_4799), .Y (n_4800));
AOI21X1 g38256(.A0 (u6_mem_b1_b_88 ), .A1 (n_5112), .B0 (n_2697), .Y(n_5054));
AOI21X1 g38251(.A0 (u7_mem_b3_b_140 ), .A1 (n_5145), .B0 (n_3242), .Y(n_5057));
AOI21X1 g38250(.A0 (u8_mem_b1_b_71 ), .A1 (n_4387), .B0 (n_2028), .Y(n_4388));
XOR2X1 g37205(.A (n_1424), .B (n_4795), .Y (n_4796));
AOI21X1 g38252(.A0 (u6_mem_b3_b_146 ), .A1 (n_5100), .B0 (n_3180), .Y(n_5056));
NAND2X1 g37759(.A (n_3215), .B (n_3214), .Y (n_4589));
NAND2X1 g37758(.A (n_3536), .B (n_2312), .Y (n_4590));
AOI21X1 g37209(.A0 (n_5526), .A1 (n_6649), .B0 (n_4675), .Y (n_5527));
MX2X1 g37208(.A (u11_mem_b1_b_149 ), .B (n_5300), .S0 (n_6502), .Y(n_5381));
AOI21X1 g38259(.A0 (u6_mem_b3_b_143 ), .A1 (n_5059), .B0 (n_3169), .Y(n_5052));
AOI21X1 g38258(.A0 (u6_mem_b3_b_144 ), .A1 (n_5059), .B0 (n_3228), .Y(n_5053));
OAI21X1 g33040(.A0 (n_7241), .A1 (n_7089), .B0 (n_12504), .Y(n_10206));
OAI21X1 g33043(.A0 (n_12483), .A1 (n_7084), .B0 (n_12504), .Y(n_10201));
OAI21X1 g33042(.A0 (n_7239), .A1 (n_7085), .B0 (n_12161), .Y(n_10202));
OAI21X1 g33045(.A0 (n_7235), .A1 (n_7181), .B0 (n_12504), .Y(n_10199));
OAI21X1 g33044(.A0 (n_7236), .A1 (n_7182), .B0 (n_12504), .Y(n_10200));
OAI21X1 g33047(.A0 (n_7232), .A1 (n_7178), .B0 (n_12504), .Y(n_10196));
OAI21X1 g33046(.A0 (n_7233), .A1 (n_7179), .B0 (n_12504), .Y(n_10198));
NAND2X1 g39337(.A (n_12826), .B (u3_mem_b0_b_101 ), .Y (n_11721));
INVX1 g42165(.A (u11_mem_b1_b ), .Y (n_6522));
NOR2X1 g39336(.A (n_3089), .B (n_2763), .Y (n_3865));
MX2X1 g36170(.A (n_5951), .B (n_5987), .S0 (n_6359), .Y (n_5952));
CLKBUFX3 g45499(.A (n_552), .Y (n_12076));
AOI21X1 g38205(.A0 (u8_mem_b1_b_62 ), .A1 (n_4502), .B0 (n_2058), .Y(n_4402));
AND2X1 g37513(.A (n_1262), .B (n_1284), .Y (n_1285));
NOR2X1 g40186(.A (n_2054), .B (n_2732), .Y (n_2055));
NOR2X1 g40187(.A (n_2684), .B (n_2118), .Y (n_2053));
NOR2X1 g40184(.A (n_2720), .B (n_1985), .Y (n_2056));
NOR2X1 g40185(.A (n_2788), .B (n_2748), .Y (n_2728));
NOR2X1 g40182(.A (n_2784), .B (n_2686), .Y (n_2731));
NOR2X1 g40183(.A (n_2751), .B (n_2729), .Y (n_2730));
NOR2X1 g40180(.A (n_2804), .B (n_2057), .Y (n_2058));
NOR2X1 g40181(.A (n_1226), .B (n_2732), .Y (n_2734));
NOR2X1 g40188(.A (n_1147), .B (n_2765), .Y (n_2727));
NOR2X1 g40189(.A (n_2477), .B (n_2748), .Y (n_1632));
NAND2X1 g36994(.A (n_1567), .B (n_1566), .Y (n_4001));
NAND2X1 g41581(.A (u26_ps_cnt_b3_b ), .B (n_760), .Y (n_910));
OR2X1 g41580(.A (n_11762), .B (n_1119), .Y (n_1120));
NOR2X1 g41582(.A (u13_ints_r_b7_b ), .B (n_488), .Y (n_550));
NOR2X1 g37512(.A (n_4764), .B (n_5371), .Y (n_3955));
MX2X1 g36150(.A (n_6392), .B (n_6533), .S0 (n_6856), .Y (n_6393));
MX2X1 g36151(.A (n_6390), .B (n_6586), .S0 (n_6341), .Y (n_6391));
MX2X1 g36152(.A (n_6388), .B (n_6453), .S0 (n_6359), .Y (n_6389));
MX2X1 g36153(.A (n_5962), .B (n_6017), .S0 (n_6341), .Y (n_5963));
MX2X1 g36154(.A (n_5959), .B (n_5997), .S0 (n_6341), .Y (n_5960));
MX2X1 g36155(.A (n_6386), .B (n_6602), .S0 (n_6341), .Y (n_6387));
MX2X1 g36156(.A (n_6384), .B (n_6599), .S0 (n_6341), .Y (n_6385));
MX2X1 g36157(.A (n_6382), .B (n_6596), .S0 (n_6341), .Y (n_6383));
MX2X1 g36158(.A (n_6380), .B (n_6592), .S0 (n_6341), .Y (n_6381));
MX2X1 g36159(.A (n_6377), .B (n_6521), .S0 (n_6359), .Y (n_6378));
NAND2X1 g36404(.A (n_5707), .B (n_6318), .Y (n_6271));
NAND2X1 g36403(.A (n_5898), .B (n_2567), .Y (n_5905));
NAND2X1 g36400(.A (n_6159), .B (n_2567), .Y (n_6275));
NAND2X1 g36401(.A (n_6204), .B (n_12634), .Y (n_12046));
NAND2X1 g39072(.A (n_12369), .B (u6_mem_b0_b_118 ), .Y (n_3472));
INVX1 g42726(.A (n_991), .Y (n_5831));
INVX2 g42727(.A (n_2343), .Y (n_10940));
INVX2 g42721(.A (oc0_cfg), .Y (n_459));
INVX1 g31759(.A (n_10341), .Y (n_10794));
AOI21X1 g31758(.A0 (n_9620), .A1 (i4_full), .B0 (n_608), .Y (n_9968));
NAND2X1 g40989(.A (n_487), .B (u11_wp_b1_b ), .Y (n_1157));
INVX1 g31753(.A (n_10795), .Y (n_10904));
NAND3X1 g31752(.A (n_6773), .B (n_12503), .C (n_1481), .Y (n_11105));
AOI21X1 g31751(.A0 (n_9534), .A1 (n_12161), .B0 (n_668), .Y(n_10796));
INVX1 g31750(.A (n_10796), .Y (n_10905));
INVX1 g31757(.A (n_9968), .Y (n_10342));
AOI21X1 g31756(.A0 (i3_full), .A1 (n_9690), .B0 (n_739), .Y (n_9694));
INVX1 g31755(.A (n_9694), .Y (n_9758));
AOI21X1 g31754(.A0 (n_9532), .A1 (n_10483), .B0 (n_611), .Y(n_10795));
AOI21X1 g30808(.A0 (n_12006), .A1 (n_12007), .B0 (n_1473), .Y(n_10928));
AND2X1 g30809(.A (n_9964), .B (n_11600), .Y (n_10801));
NOR2X1 g35838(.A (n_5632), .B (n_1777), .Y (n_5624));
XOR2X1 g40401(.A (n_6838), .B (n_814), .Y (n_1833));
NOR2X1 g41639(.A (u2_res_cnt_b1_b ), .B (u2_res_cnt_b3_b ), .Y (n_415));
AOI21X1 g30800(.A0 (n_12012), .A1 (n_12013), .B0 (n_1473), .Y(n_10934));
NOR2X1 g30801(.A (n_10791), .B (n_10940), .Y (n_10999));
NOR2X1 g30802(.A (n_10789), .B (n_10940), .Y (n_10998));
AOI21X1 g30803(.A0 (n_12140), .A1 (n_11536), .B0 (n_1473), .Y(n_10933));
AOI21X1 g30804(.A0 (n_12150), .A1 (n_11538), .B0 (n_10940), .Y(n_10932));
AOI21X1 g30805(.A0 (n_12042), .A1 (n_12043), .B0 (n_10940), .Y(n_10931));
AOI21X1 g30806(.A0 (n_11950), .A1 (n_11951), .B0 (n_10945), .Y(n_10930));
AOI21X1 g30807(.A0 (n_11980), .A1 (n_11981), .B0 (n_1473), .Y(n_10929));
NAND2X1 g37540(.A (n_620), .B (in_slt_742), .Y (n_1010));
NAND2X1 g37541(.A (n_531), .B (in_slt_742), .Y (n_1009));
INVX1 g43002(.A (u11_mem_b1_b_124 ), .Y (n_6487));
NOR2X1 g37542(.A (n_4743), .B (n_5371), .Y (n_3952));
NAND2X1 g39070(.A (u6_mem_b2_b_47 ), .B (n_3474), .Y (n_12818));
INVX1 g43003(.A (u14_n_134), .Y (n_1124));
INVX1 g42588(.A (u11_mem_b0_b_171 ), .Y (n_1755));
NOR2X1 g40964(.A (n_1924), .B (n_1424), .Y (n_1425));
INVX8 g40965(.A (n_1158), .Y (n_6898));
NAND2X1 g37544(.A (n_539), .B (in_slt_742), .Y (n_1008));
INVX1 g43001(.A (u9_mem_b2_b ), .Y (n_509));
INVX1 g42585(.A (u10_mem_b1_b_130 ), .Y (n_6463));
INVX1 g42586(.A (u11_mem_b3_b_83 ), .Y (n_5502));
NAND4X1 g37097(.A (n_11453), .B (n_11454), .C (n_3374), .D (n_2391),.Y (n_6182));
NAND2X1 g37546(.A (n_5480), .B (n_3492), .Y (n_4646));
NAND2X1 g37547(.A (n_843), .B (in_slt_742), .Y (n_1260));
AOI21X1 g38236(.A0 (u6_mem_b3_b_152 ), .A1 (n_5059), .B0 (n_3022), .Y(n_5063));
NOR2X1 g40263(.A (n_2721), .B (n_2691), .Y (n_2692));
NOR2X1 g41164(.A (n_1198), .B (u8_wp_b0_b ), .Y (n_920));
NOR2X1 g40262(.A (n_938), .B (n_2707), .Y (n_2001));
NAND2X2 g41163(.A (n_473), .B (n_751), .Y (n_1147));
AOI22X1 g37658(.A0 (u9_din_tmp_55), .A1 (n_2368), .B0 (in_slt_410),.B1 (n_3935), .Y (n_3934));
NOR2X1 g39122(.A (n_2831), .B (n_1488), .Y (n_1498));
INVX2 g41162(.A (n_1147), .Y (n_1409));
NAND2X1 g39577(.A (u5_mem_b1_b_86 ), .B (n_3239), .Y (n_3087));
NAND2X1 g39576(.A (n_2330), .B (u7_mem_b0_b_100 ), .Y (n_2281));
NAND2X1 g39575(.A (u6_mem_b2_b_39 ), .B (n_2285), .Y (n_2282));
NAND2X1 g39573(.A (u6_mem_b1_b_70 ), .B (n_12169), .Y (n_11708));
INVX4 g39571(.A (n_2284), .Y (n_5591));
NOR2X1 g40267(.A (n_2470), .B (n_3008), .Y (n_1999));
AOI21X1 g38185(.A0 (u4_mem_b3_b_131 ), .A1 (n_5106), .B0 (n_2882), .Y(n_5107));
NAND2X1 g39578(.A (u6_mem_b1_b_83 ), .B (n_4253), .Y (n_4165));
MX2X1 g34127(.A (u8_mem_b0_b_102 ), .B (n_3817), .S0 (n_7490), .Y(n_9383));
MX2X1 g34126(.A (u8_mem_b0_b_101 ), .B (n_3814), .S0 (n_7490), .Y(n_9385));
MX2X1 g34125(.A (u3_mem_b0_b_107 ), .B (n_3815), .S0 (n_8700), .Y(n_8720));
MX2X1 g34124(.A (u8_mem_b0_b_100 ), .B (n_3602), .S0 (n_7490), .Y(n_8721));
MX2X1 g34123(.A (u8_mem_b0_b ), .B (n_3604), .S0 (n_7490), .Y(n_9386));
MX2X1 g34122(.A (u3_mem_b0_b_106 ), .B (n_3603), .S0 (n_7423), .Y(n_8722));
MX2X1 g34121(.A (u3_mem_b0_b_105 ), .B (n_3804), .S0 (n_8700), .Y(n_9387));
MX2X1 g34120(.A (u3_mem_b0_b_104 ), .B (n_3813), .S0 (n_7423), .Y(n_8252));
AOI22X1 g37659(.A0 (u9_din_tmp_56), .A1 (n_2368), .B0 (in_slt_411),.B1 (n_3935), .Y (n_3933));
INVX1 g41617(.A (n_977), .Y (n_1116));
MX2X1 g34129(.A (u8_mem_b0_b_103 ), .B (n_3818), .S0 (n_7490), .Y(n_8718));
MX2X1 g34128(.A (u3_mem_b0_b_108 ), .B (n_3601), .S0 (n_8700), .Y(n_8719));
NAND2X1 g34390(.A (u4_mem_b2_b_41 ), .B (n_7984), .Y (n_8014));
OAI21X1 g33656(.A0 (n_4359), .A1 (n_9212), .B0 (n_7884), .Y (n_9250));
NAND2X1 g39074(.A (in_slt_407), .B (n_2368), .Y (n_4757));
NAND2X1 g34391(.A (u4_mem_b2_b_42 ), .B (n_7984), .Y (n_8013));
NOR2X1 g35854(.A (n_4087), .B (n_5442), .Y (n_5443));
NAND2X1 g34392(.A (u4_mem_b2_b_43 ), .B (n_7984), .Y (n_8012));
NAND2X1 g34393(.A (n_6681), .B (n_7462), .Y (n_8228));
OAI21X1 g35857(.A0 (n_2615), .A1 (u2_to_cnt_b5_b ), .B0 (n_2616), .Y(n_4853));
NAND2X1 g34395(.A (u4_mem_b2_b_45 ), .B (n_7984), .Y (n_8010));
NOR2X1 g39753(.A (n_3332), .B (n_2712), .Y (n_2977));
AOI21X1 g35674(.A0 (i4_dout_622), .A1 (n_7468), .B0 (n_7108), .Y(n_7299));
NAND2X1 g39751(.A (n_3339), .B (in_slt_431), .Y (n_5355));
INVX1 g39750(.A (n_5355), .Y (n_4135));
NAND2X1 g39757(.A (n_11789), .B (u8_mem_b0_b_119 ), .Y (n_2974));
NAND2X1 g34396(.A (u4_mem_b2_b_46 ), .B (n_7984), .Y (n_8009));
NAND2X1 g39755(.A (u8_mem_b2_b_45 ), .B (n_2362), .Y (n_2253));
OAI21X1 g35859(.A0 (n_5728), .A1 (n_11934), .B0 (n_6815), .Y(n_7202));
MX2X1 g38668(.A (u5_mem_b0_b_121 ), .B (wb_din_691), .S0 (n_3720), .Y(n_3698));
NAND2X1 g39759(.A (n_2325), .B (in_slt_444), .Y (n_2251));
NAND2X1 g34465(.A (u4_mem_b3_b_124 ), .B (n_7984), .Y (n_7956));
MX2X1 g38669(.A (u5_mem_b0_b_93 ), .B (wb_din_663), .S0 (n_3720), .Y(n_3697));
OAI21X1 g33863(.A0 (n_4541), .A1 (n_9034), .B0 (n_7663), .Y (n_8992));
OAI21X1 g33862(.A0 (n_4538), .A1 (n_9034), .B0 (n_7664), .Y (n_8993));
OAI21X1 g33861(.A0 (n_4536), .A1 (n_9010), .B0 (n_8145), .Y (n_8995));
OAI21X1 g33860(.A0 (n_4309), .A1 (n_9043), .B0 (n_7665), .Y (n_8996));
OAI21X1 g33867(.A0 (n_4366), .A1 (n_8948), .B0 (n_7658), .Y (n_8988));
OAI21X1 g33866(.A0 (n_4339), .A1 (n_9043), .B0 (n_7659), .Y (n_8989));
OAI21X1 g33865(.A0 (n_4546), .A1 (n_9034), .B0 (n_7660), .Y (n_8990));
OAI21X1 g33864(.A0 (n_4307), .A1 (n_8981), .B0 (n_7661), .Y (n_8991));
AOI21X1 g35670(.A0 (i3_dout_587), .A1 (n_6700), .B0 (n_7110), .Y(n_7303));
OAI21X1 g33869(.A0 (n_4292), .A1 (n_9010), .B0 (n_7656), .Y (n_8986));
OAI21X1 g33868(.A0 (n_4305), .A1 (n_8948), .B0 (n_7657), .Y (n_8987));
AOI21X1 g35671(.A0 (i3_dout_588), .A1 (n_6700), .B0 (n_7106), .Y(n_7386));
MX2X1 g38664(.A (u5_mem_b0_b_118 ), .B (wb_din_688), .S0 (n_3720), .Y(n_3707));
AOI21X1 g35672(.A0 (i4_dout_620), .A1 (n_7468), .B0 (n_7045), .Y(n_7301));
MX2X1 g38665(.A (u5_mem_b0_b_119 ), .B (wb_din_689), .S0 (n_841), .Y(n_3704));
AOI21X1 g35673(.A0 (i4_dout_621), .A1 (n_7468), .B0 (n_7109), .Y(n_7300));
MX2X1 g38666(.A (u5_mem_b0_b_92 ), .B (wb_din_662), .S0 (n_841), .Y(n_3700));
INVX1 g42167(.A (u11_mem_b2_b_89 ), .Y (n_6448));
MX2X1 g38667(.A (u5_mem_b0_b_120 ), .B (wb_din_690), .S0 (n_3720), .Y(n_3699));
NAND2X1 g37654(.A (n_2459), .B (n_2636), .Y (n_4627));
NAND2X1 g37140(.A (n_4621), .B (n_3351), .Y (n_6920));
MX2X1 g38661(.A (u5_mem_b0_b_115 ), .B (wb_din_685), .S0 (n_841), .Y(n_3712));
MX2X1 g38662(.A (u7_mem_b0_b ), .B (wb_din), .S0 (n_3622), .Y(n_3710));
MX2X1 g38663(.A (u5_mem_b0_b_116 ), .B (wb_din_686), .S0 (n_3720), .Y(n_3709));
AOI22X1 g37324(.A0 (n_4729), .A1 (oc4_cfg_1004), .B0 (n_5591), .B1(ic0_cfg_1024), .Y (n_4730));
AOI22X1 g37655(.A0 (n_2558), .A1 (n_5959), .B0 (n_5998), .B1(n_2544), .Y (n_1862));
AOI21X1 g38517(.A0 (u7_mem_b3_b_144 ), .A1 (n_4961), .B0 (n_3324), .Y(n_4882));
AOI22X1 g37326(.A0 (n_5277), .A1 (crac_out_865), .B0 (n_6972), .B1(oc2_cfg_987), .Y (n_4728));
AOI22X1 g37327(.A0 (n_5272), .A1 (u13_intm_r_b20_b ), .B0(u13_ints_r_b20_b ), .B1 (n_4726), .Y (n_4727));
NAND2X1 g37896(.A (n_4236), .B (n_3104), .Y (n_5196));
AOI21X1 g38119(.A0 (u7_mem_b1_b_61 ), .A1 (n_5118), .B0 (n_2783), .Y(n_5119));
AOI21X1 g38513(.A0 (u8_mem_b1_b_66 ), .A1 (n_4387), .B0 (n_2046), .Y(n_4302));
NOR2X1 g40216(.A (n_938), .B (n_2831), .Y (n_2034));
NOR2X1 g40217(.A (n_945), .B (n_2772), .Y (n_2032));
NOR2X1 g40214(.A (n_2713), .B (n_2712), .Y (n_2714));
NOR2X1 g40215(.A (n_2103), .B (n_2744), .Y (n_2035));
NOR2X1 g40212(.A (n_2792), .B (n_933), .Y (n_2036));
AOI22X1 g37322(.A0 (n_5272), .A1 (u13_intm_r_b17_b ), .B0(u13_ints_r_b17_b ), .B1 (n_4726), .Y (n_4731));
NOR2X1 g40210(.A (n_2038), .B (n_2767), .Y (n_2039));
NOR2X1 g40211(.A (n_2081), .B (n_2765), .Y (n_2037));
AOI21X1 g38511(.A0 (u7_mem_b3_b_135 ), .A1 (n_5145), .B0 (n_2930), .Y(n_4886));
AOI22X1 g37751(.A0 (n_2558), .A1 (n_1238), .B0 (n_5352), .B1(n_1316), .Y (n_1239));
NOR2X1 g40219(.A (n_1226), .B (n_2702), .Y (n_2711));
INVX2 g40624(.A (wb_din_686), .Y (n_2702));
NAND2X1 g39951(.A (n_12369), .B (u6_mem_b0_b_93 ), .Y (n_2855));
NAND2X1 g34378(.A (u4_mem_b1_b_62 ), .B (n_7984), .Y (n_8025));
NOR2X1 g39953(.A (n_3117), .B (n_2772), .Y (n_2854));
NAND2X1 g38849(.A (u5_mem_b3_b_147 ), .B (n_3543), .Y (n_2443));
NAND4X1 g45932(.A (n_12674), .B (n_12675), .C (n_12676), .D(n_12680), .Y (n_12681));
NAND2X1 g39952(.A (u6_mem_b2_b ), .B (n_2285), .Y (n_2229));
NAND2X1 g45934(.A (n_12823), .B (u5_mem_b2_b_46 ), .Y (n_12675));
NAND2X1 g45936(.A (n_12679), .B (u5_mem_b0_b_108 ), .Y (n_12680));
CLKBUFX3 g45937(.A (n_12678), .Y (n_12679));
INVX2 g45938(.A (n_12677), .Y (n_12678));
NOR2X1 g39955(.A (n_2702), .B (n_1488), .Y (n_1555));
AOI22X1 g37650(.A0 (n_6902), .A1 (n_1835), .B0 (n_6912), .B1(n_1760), .Y (n_1710));
NAND2X1 g39954(.A (n_11798), .B (u8_mem_b0_b_101 ), .Y (n_11459));
NOR2X1 g40378(.A (n_1226), .B (n_2864), .Y (n_2647));
NOR2X1 g40375(.A (n_2794), .B (n_2045), .Y (n_1930));
NOR2X1 g40374(.A (n_2792), .B (n_1985), .Y (n_1931));
NOR2X1 g40377(.A (n_1016), .B (n_2691), .Y (n_2648));
NAND2X1 g39956(.A (u8_mem_b1_b_83 ), .B (n_12291), .Y (n_2852));
NOR2X1 g40371(.A (n_2085), .B (n_2786), .Y (n_1934));
NOR2X1 g40370(.A (n_2006), .B (n_2691), .Y (n_1935));
NOR2X1 g40373(.A (n_2171), .B (n_2818), .Y (n_1932));
NOR2X1 g40372(.A (n_2054), .B (n_2755), .Y (n_1933));
AOI21X1 g38008(.A0 (u3_mem_b1_b_66 ), .A1 (n_5157), .B0 (n_2651), .Y(n_5150));
AOI21X1 g38009(.A0 (u3_mem_b1_b_67 ), .A1 (n_5148), .B0 (n_2781), .Y(n_5149));
AOI21X1 g38000(.A0 (u8_mem_b3_b_134 ), .A1 (n_3879), .B0 (n_1458), .Y(n_3889));
AOI21X1 g38001(.A0 (u3_mem_b1_b_62 ), .A1 (n_5157), .B0 (n_2789), .Y(n_5154));
AOI21X1 g38002(.A0 (u3_mem_b1_b_63 ), .A1 (n_5157), .B0 (n_2718), .Y(n_5153));
AOI21X1 g38003(.A0 (u7_mem_b2_b_58 ), .A1 (n_4540), .B0 (n_2222), .Y(n_4541));
AOI21X1 g38004(.A0 (u3_mem_b1_b_64 ), .A1 (n_5148), .B0 (n_2679), .Y(n_5152));
AOI21X1 g38005(.A0 (u6_mem_b2_b_52 ), .A1 (n_4544), .B0 (n_2219), .Y(n_4539));
AOI21X1 g38006(.A0 (u3_mem_b1_b_65 ), .A1 (n_5157), .B0 (n_2776), .Y(n_5151));
AOI21X1 g38007(.A0 (u8_mem_b3_b_141 ), .A1 (n_3879), .B0 (n_1504), .Y(n_3888));
NAND2X1 g37752(.A (n_3528), .B (n_2235), .Y (n_4593));
AND2X1 g45463(.A (n_634), .B (n_12535), .Y (n_11912));
AND2X1 g30789(.A (n_10340), .B (n_11772), .Y (n_10948));
AOI22X1 g37755(.A0 (n_196), .A1 (n_2530), .B0 (n_2542), .B1 (n_2534),.Y (n_2543));
AOI22X1 g37653(.A0 (n_6893), .A1 (n_1835), .B0 (n_6905), .B1(n_1760), .Y (n_1706));
AOI22X1 g37754(.A0 (n_6884), .A1 (n_1859), .B0 (n_6873), .B1(n_1835), .Y (n_1836));
INVX2 g36903(.A (n_5713), .Y (n_5714));
NAND2X1 g39130(.A (u8_mem_b2_b_38 ), .B (n_2362), .Y (n_2353));
NAND2X1 g36366(.A (n_6814), .B (n_6824), .Y (n_6819));
OAI21X1 g33788(.A0 (n_5006), .A1 (n_9087), .B0 (n_7739), .Y (n_9086));
OAI21X1 g33789(.A0 (n_5061), .A1 (n_9087), .B0 (n_7738), .Y (n_9085));
NAND2X1 g36363(.A (n_6167), .B (n_6316), .Y (n_6304));
NAND2X1 g36362(.A (n_5837), .B (n_6821), .Y (n_5917));
NAND2X1 g36361(.A (n_5841), .B (n_6821), .Y (n_5918));
NAND2X1 g36360(.A (n_5544), .B (n_12634), .Y (n_5919));
OAI21X1 g33782(.A0 (n_5052), .A1 (n_9165), .B0 (n_7745), .Y (n_9094));
OAI21X1 g33783(.A0 (n_5053), .A1 (n_9165), .B0 (n_7744), .Y (n_9093));
OAI21X1 g33780(.A0 (n_5051), .A1 (n_9165), .B0 (n_7747), .Y (n_9097));
OAI21X1 g33781(.A0 (n_4921), .A1 (n_9165), .B0 (n_7746), .Y (n_9096));
OAI21X1 g33786(.A0 (n_4920), .A1 (n_9087), .B0 (n_7741), .Y (n_9089));
NAND2X1 g34372(.A (u4_mem_b1_b_87 ), .B (n_7984), .Y (n_8030));
OAI21X1 g33784(.A0 (n_5055), .A1 (n_9105), .B0 (n_7743), .Y (n_9092));
OAI21X1 g33785(.A0 (n_5056), .A1 (n_9105), .B0 (n_7742), .Y (n_9091));
MX2X1 g31322(.A (n_5659), .B (n_1581), .S0 (n_10513), .Y (n_10428));
MX2X1 g31323(.A (n_5646), .B (n_2550), .S0 (n_9724), .Y (n_10426));
MX2X1 g31320(.A (n_5647), .B (n_1685), .S0 (n_10137), .Y (n_10128));
MX2X1 g31321(.A (n_5648), .B (n_1585), .S0 (n_10513), .Y (n_10429));
MX2X1 g31326(.A (n_5471), .B (n_1677), .S0 (n_9724), .Y (n_10423));
XOR2X1 g31327(.A (n_784), .B (n_9902), .Y (n_10811));
MX2X1 g31324(.A (n_6356), .B (n_6355), .S0 (n_10513), .Y (n_10425));
MX2X1 g31325(.A (n_6354), .B (n_6353), .S0 (n_10513), .Y (n_10424));
MX2X1 g31328(.A (n_6352), .B (n_6351), .S0 (n_10537), .Y (n_10422));
MX2X1 g31329(.A (n_5470), .B (n_1240), .S0 (n_9724), .Y (n_10421));
NAND2X1 g37944(.A (n_3548), .B (n_3399), .Y (n_12852));
NAND2X1 g37945(.A (n_3499), .B (n_3482), .Y (n_5191));
INVX1 g37414(.A (n_3943), .Y (n_4680));
INVX1 g37415(.A (n_4634), .Y (n_5250));
OAI21X1 g37412(.A0 (u9_mem_b0_b_171 ), .A1 (n_6856), .B0 (n_4639), .Y(n_5468));
NAND2X1 g37941(.A (n_3354), .B (n_2957), .Y (n_5193));
OAI21X1 g37410(.A0 (u10_mem_b0_b_180 ), .A1 (n_6341), .B0 (n_5228), .Y(n_5641));
OAI21X1 g37411(.A0 (u10_mem_b0_b_178 ), .A1 (n_6341), .B0 (n_5229), .Y(n_5639));
NAND2X1 g37948(.A (n_2437), .B (n_3331), .Y (n_5190));
NAND2X1 g37949(.A (n_2389), .B (n_2367), .Y (n_4553));
XOR2X1 g37418(.A (n_6838), .B (n_763), .Y (n_1269));
XOR2X1 g37419(.A (n_614), .B (n_765), .Y (n_1790));
CLKBUFX3 g41134(.A (n_1149), .Y (n_2285));
INVX1 g41130(.A (n_969), .Y (n_1045));
CLKBUFX1 g41132(.A (n_969), .Y (n_5730));
NOR2X1 g41133(.A (n_689), .B (u9_wp_b2_b ), .Y (n_969));
INVX2 g41138(.A (n_1411), .Y (n_3474));
MX2X1 g36090(.A (n_6490), .B (n_6442), .S0 (n_6502), .Y (n_6491));
MX2X1 g36093(.A (n_5984), .B (n_5983), .S0 (n_6502), .Y (n_5985));
MX2X1 g36092(.A (n_6484), .B (n_6483), .S0 (n_6502), .Y (n_6485));
MX2X1 g36095(.A (n_419), .B (n_6521), .S0 (n_5312), .Y (n_6481));
MX2X1 g36094(.A (n_5981), .B (n_5997), .S0 (n_6475), .Y (n_5982));
MX2X1 g36097(.A (n_6476), .B (n_6602), .S0 (n_6475), .Y (n_6477));
MX2X1 g36096(.A (n_6479), .B (n_6478), .S0 (n_5312), .Y (n_6480));
MX2X1 g36099(.A (n_6471), .B (n_6514), .S0 (n_5409), .Y (n_6472));
MX2X1 g36098(.A (n_433), .B (n_6473), .S0 (n_5312), .Y (n_6474));
INVX1 g39772(.A (n_4751), .Y (n_2968));
AOI22X1 g37892(.A0 (u11_din_tmp_55), .A1 (n_4560), .B0 (n_4097), .B1(in_slt_456), .Y (n_3900));
AOI22X1 g37893(.A0 (u10_din_tmp_55), .A1 (n_3339), .B0 (n_3911), .B1(in_slt_434), .Y (n_3899));
AOI22X1 g37365(.A0 (n_5272), .A1 (u13_intm_r_b15_b ), .B0 (n_5277),.B1 (crac_din_706), .Y (n_5253));
AOI21X1 g38346(.A0 (u7_mem_b1_b_79 ), .A1 (n_5118), .B0 (n_2734), .Y(n_4991));
AOI22X1 g37890(.A0 (n_2558), .A1 (n_6342), .B0 (n_6578), .B1(n_1316), .Y (n_1295));
INVX1 g42112(.A (u9_mem_b3_b_77 ), .Y (n_5374));
INVX1 g42111(.A (oc0_cfg_966), .Y (n_925));
NAND2X1 g34808(.A (u7_mem_b3_b_125 ), .B (n_7651), .Y (n_7625));
NAND2X1 g34809(.A (u7_mem_b3_b_126 ), .B (n_7651), .Y (n_7624));
INVX1 g42115(.A (u10_mem_b0_b_162 ), .Y (n_6380));
NAND2X1 g34804(.A (u8_mem_b3_b_137 ), .B (n_7976), .Y (n_7629));
NAND2X1 g34805(.A (u7_mem_b3_b_151 ), .B (n_7651), .Y (n_7628));
NAND2X1 g34806(.A (u7_mem_b3_b_152 ), .B (n_7651), .Y (n_7627));
NAND2X1 g34807(.A (u7_mem_b3_b_124 ), .B (n_7651), .Y (n_7626));
NAND2X1 g34800(.A (u7_mem_b3_b_148 ), .B (n_7651), .Y (n_7633));
NAND2X1 g34801(.A (u7_mem_b3_b_149 ), .B (n_7651), .Y (n_7632));
NAND2X1 g34802(.A (u7_mem_b3_b_150 ), .B (n_7651), .Y (n_7631));
NAND2X1 g34803(.A (u7_mem_b3_b_123 ), .B (n_7651), .Y (n_7630));
NOR2X1 g35318(.A (in_valid_s_b0_b ), .B (n_1308), .Y (n_9352));
OR2X1 g35317(.A (n_11827), .B (n_12585), .Y (n_8660));
NOR2X1 g35316(.A (n_7017), .B (n_12335), .Y (n_7537));
INVX1 g35315(.A (n_7537), .Y (n_8661));
INVX1 g35314(.A (n_8661), .Y (n_9475));
OR2X1 g35313(.A (n_5825), .B (n_11827), .Y (n_8662));
NOR2X1 g35312(.A (n_1100), .B (n_12335), .Y (n_7538));
INVX1 g35311(.A (n_7538), .Y (n_8663));
INVX1 g35310(.A (n_8663), .Y (n_9476));
NAND2X1 g36958(.A (n_2563), .B (n_3930), .Y (n_5382));
NAND2X1 g36959(.A (n_1593), .B (n_1590), .Y (n_4010));
NAND2X1 g36950(.A (n_1616), .B (n_1613), .Y (n_4015));
NAND2X1 g36951(.A (n_1611), .B (n_1607), .Y (n_4014));
NAND2X1 g36952(.A (n_2525), .B (n_2523), .Y (n_4808));
NAND2X1 g36953(.A (n_1606), .B (n_1603), .Y (n_4013));
NAND2X1 g36954(.A (n_1601), .B (n_1855), .Y (n_4012));
INVX1 g36955(.A (n_6161), .Y (n_5705));
NAND4X1 g36956(.A (n_2927), .B (n_2924), .C (n_3143), .D (n_2402), .Y(n_6161));
NAND2X1 g36957(.A (n_1597), .B (n_1594), .Y (n_4011));
AOI22X1 g37897(.A0 (n_4097), .A1 (in_slt_459), .B0 (n_2325), .B1(in_slt_457), .Y (n_2516));
AOI21X1 g38342(.A0 (u5_mem_b3_b_135 ), .A1 (n_4996), .B0 (n_2934), .Y(n_4995));
AOI22X1 g37894(.A0 (n_3911), .A1 (in_slt_437), .B0 (n_2344), .B1(in_slt_435), .Y (n_2519));
NAND2X1 g26(.A (n_4829), .B (n_2568), .Y (n_12588));
INVX2 g24(.A (valid_s), .Y (n_12335));
NOR2X1 g25(.A (n_12589), .B (n_10663), .Y (n_12590));
INVX1 g22(.A (n_12336), .Y (n_12340));
NOR2X1 g23(.A (n_11128), .B (n_12591), .Y (n_12592));
INVX1 g20(.A (dma_ack_i_b6_b), .Y (n_12370));
NAND4X1 g28(.A (n_12361), .B (n_12362), .C (n_12363), .D (n_12367),.Y (n_12368));
AOI22X1 g29(.A0 (u4_mem_b3_b_136 ), .A1 (n_12744), .B0 (n_12273), .B1(u4_mem_b1_b_74 ), .Y (n_11846));
INVX1 g42913(.A (u9_mem_b0_b_165 ), .Y (n_6866));
AOI22X1 g37895(.A0 (n_4097), .A1 (in_slt_458), .B0 (n_2325), .B1(in_slt_456), .Y (n_2517));
NAND2X1 g34853(.A (u3_mem_b1_b_77 ), .B (n_8141), .Y (n_7581));
OAI21X1 g33418(.A0 (n_3847), .A1 (n_8453), .B0 (n_7629), .Y (n_8454));
OAI21X1 g33419(.A0 (n_5152), .A1 (n_8097), .B0 (n_8158), .Y (n_8452));
OAI21X1 g33412(.A0 (n_3842), .A1 (n_8930), .B0 (n_7609), .Y (n_8462));
OAI21X1 g33413(.A0 (n_5154), .A1 (n_8911), .B0 (n_8164), .Y (n_8460));
NAND2X1 g34370(.A (u4_mem_b1_b_85 ), .B (n_7984), .Y (n_8032));
OAI21X1 g33411(.A0 (n_5155), .A1 (n_8856), .B0 (n_7607), .Y (n_8463));
NAND2X1 g34376(.A (u4_mem_b1_b_90 ), .B (n_7984), .Y (n_8026));
NAND2X1 g34377(.A (n_6684), .B (n_7464), .Y (n_8230));
OAI21X1 g33414(.A0 (n_3889), .A1 (n_8457), .B0 (n_8163), .Y (n_8459));
NAND2X1 g34375(.A (u4_mem_b1_b_89 ), .B (n_7984), .Y (n_8027));
AOI21X1 g38493(.A0 (u7_mem_b2_b_41 ), .A1 (n_4509), .B0 (n_1995), .Y(n_4317));
AOI21X1 g38492(.A0 (u7_mem_b2_b_39 ), .A1 (n_4540), .B0 (n_2064), .Y(n_4318));
AOI21X1 g38491(.A0 (u7_mem_b1_b_68 ), .A1 (n_5118), .B0 (n_2688), .Y(n_4890));
AOI21X1 g38490(.A0 (u8_mem_b1_b_87 ), .A1 (n_4502), .B0 (n_1946), .Y(n_4319));
AOI21X1 g38495(.A0 (u3_mem_b3_b_133 ), .A1 (n_5133), .B0 (n_2912), .Y(n_4889));
AOI21X1 g38494(.A0 (u7_mem_b2_b_42 ), .A1 (n_4509), .B0 (n_2060), .Y(n_4316));
AOI21X1 g38499(.A0 (u7_mem_b2_b_53 ), .A1 (n_4509), .B0 (n_2034), .Y(n_4312));
AOI21X1 g38498(.A0 (u7_mem_b2_b_47 ), .A1 (n_4509), .B0 (n_1944), .Y(n_4313));
AOI21X1 g38144(.A0 (u4_mem_b2_b_38 ), .A1 (n_4439), .B0 (n_1947), .Y(n_4441));
MX2X1 g33118(.A (n_4687), .B (wb_din_674), .S0 (n_8611), .Y (n_8613));
NAND2X1 g17(.A (n_12066), .B (n_12370), .Y (n_12371));
NAND4X1 g45509(.A (n_3317), .B (n_2914), .C (n_3396), .D (n_2467), .Y(n_12111));
NAND2X1 g37778(.A (n_3537), .B (n_2897), .Y (n_4586));
AOI21X1 g38279(.A0 (u5_mem_b1_b_79 ), .A1 (n_5037), .B0 (n_2778), .Y(n_5032));
AOI21X1 g32708(.A0 (n_6265), .A1 (n_6229), .B0 (n_10617), .Y(n_10613));
AOI21X1 g38277(.A0 (u5_mem_b1_b_60 ), .A1 (n_5037), .B0 (n_2661), .Y(n_5033));
AOI21X1 g38276(.A0 (u5_mem_b1_b_78 ), .A1 (n_5037), .B0 (n_2799), .Y(n_5034));
AOI21X1 g38275(.A0 (u5_mem_b1_b_77 ), .A1 (n_5037), .B0 (n_2666), .Y(n_5035));
AOI21X1 g38274(.A0 (u6_mem_b3_b_137 ), .A1 (n_5100), .B0 (n_3296), .Y(n_5036));
AOI21X1 g38273(.A0 (u5_mem_b1_b_76 ), .A1 (n_5037), .B0 (n_2726), .Y(n_5038));
AOI21X1 g38272(.A0 (u5_mem_b1_b_75 ), .A1 (n_5048), .B0 (n_2779), .Y(n_5039));
AOI21X1 g38271(.A0 (u5_mem_b1_b_74 ), .A1 (n_5037), .B0 (n_2747), .Y(n_5040));
AOI21X1 g38270(.A0 (u6_mem_b3_b_138 ), .A1 (n_5100), .B0 (n_3357), .Y(n_5041));
OAI21X1 g33069(.A0 (n_7123), .A1 (n_7069), .B0 (n_10483), .Y(n_11619));
OAI21X1 g33068(.A0 (n_7216), .A1 (n_6983), .B0 (n_10483), .Y(n_11617));
OAI21X1 g33063(.A0 (n_7219), .A1 (n_7067), .B0 (n_10481), .Y(n_10496));
OAI21X1 g33067(.A0 (n_7121), .A1 (n_7064), .B0 (n_10483), .Y(n_11615));
OAI21X1 g33065(.A0 (n_7217), .A1 (n_7066), .B0 (n_10481), .Y(n_10493));
OAI21X1 g33064(.A0 (n_7218), .A1 (n_6984), .B0 (n_10483), .Y(n_11633));
NAND2X1 g35326(.A (n_6745), .B (n_7337), .Y (n_7476));
NAND2X1 g35327(.A (n_6718), .B (n_11564), .Y (n_7383));
AND2X1 g35324(.A (n_1230), .B (n_7030), .Y (n_11534));
NAND3X1 g35325(.A (n_7050), .B (n_5965), .C (n_2271), .Y (n_7365));
AOI21X1 g38505(.A0 (u5_mem_b2_b_32 ), .A1 (n_4370), .B0 (n_2134), .Y(n_4306));
NAND2X1 g35451(.A (n_6692), .B (n_7302), .Y (n_7450));
NAND2X1 g35320(.A (n_11600), .B (in_valid_s_b1_b ), .Y (n_7479));
NAND2X1 g39012(.A (u7_mem_b1_b_75 ), .B (n_4225), .Y (n_4247));
OR2X1 g35321(.A (n_11762), .B (n_7477), .Y (n_7478));
AOI21X1 g38143(.A0 (u4_mem_b2_b ), .A1 (n_4439), .B0 (n_2106), .Y(n_4442));
NAND2X1 g39013(.A (u8_mem_b2_b_51 ), .B (n_3441), .Y (n_2638));
NAND2X1 g39379(.A (n_12679), .B (u5_mem_b0_b_117 ), .Y (n_3224));
NAND2X1 g39378(.A (n_12840), .B (u4_mem_b0_b_113 ), .Y (n_3225));
AOI21X1 g38507(.A0 (u8_mem_b2_b_52 ), .A1 (n_4491), .B0 (n_1826), .Y(n_4304));
XOR2X1 g38432(.A (n_214), .B (n_5138), .Y (n_4333));
INVX1 g42033(.A (u11_mem_b3_b_76 ), .Y (n_5494));
AOI21X1 g38142(.A0 (u6_mem_b2_b ), .A1 (n_4544), .B0 (n_2023), .Y(n_4443));
NAND2X1 g36428(.A (n_5823), .B (n_6152), .Y (n_5890));
MX2X1 g36138(.A (n_6396), .B (n_6582), .S0 (n_6856), .Y (n_6397));
MX2X1 g36139(.A (n_6866), .B (n_6883), .S0 (n_6856), .Y (n_6867));
AOI21X1 g38438(.A0 (u6_mem_b3_b_131 ), .A1 (n_5059), .B0 (n_2916), .Y(n_4927));
NAND2X1 g36420(.A (n_6814), .B (n_12531), .Y (n_6815));
MX2X1 g36133(.A (n_6868), .B (n_6925), .S0 (n_6856), .Y (n_6869));
NAND2X1 g36422(.A (n_12746), .B (n_12531), .Y (n_6812));
MX2X1 g36131(.A (n_6406), .B (n_6563), .S0 (n_6475), .Y (n_6407));
MX2X1 g36136(.A (n_6400), .B (n_6539), .S0 (n_6856), .Y (n_6401));
MX2X1 g36137(.A (n_6398), .B (n_6637), .S0 (n_6856), .Y (n_6399));
MX2X1 g36134(.A (n_6404), .B (n_6646), .S0 (n_6856), .Y (n_6405));
NAND2X1 g36427(.A (n_6797), .B (n_12531), .Y (n_6810));
NAND2X1 g39015(.A (n_3415), .B (in_slt_405), .Y (n_3515));
INVX1 g36989(.A (n_12626), .Y (n_5550));
AND2X1 g41659(.A (n_670), .B (n_921), .Y (n_9653));
OR2X1 g41658(.A (u10_rp_b1_b ), .B (u10_rp_b0_b ), .Y (n_481));
NAND2X1 g39016(.A (n_2468), .B (n_494), .Y (n_2369));
INVX4 g41651(.A (n_673), .Y (n_1111));
NOR2X1 g41653(.A (u13_ints_r_b0_b ), .B (n_1036), .Y (n_980));
NOR2X1 g41652(.A (n_12281), .B (n_244), .Y (n_673));
INVX2 g41657(.A (n_481), .Y (n_2558));
NOR2X1 g41656(.A (n_671), .B (n_924), .Y (n_672));
INVX1 g36896(.A (n_5884), .Y (n_5563));
NAND2X1 g39017(.A (u7_mem_b2_b_46 ), .B (n_12645), .Y (n_3514));
INVX1 g39086(.A (n_5315), .Y (n_4232));
AOI21X1 g38027(.A0 (u6_mem_b2_b_48 ), .A1 (n_4544), .B0 (n_2211), .Y(n_4525));
AOI21X1 g38502(.A0 (u7_mem_b2_b_56 ), .A1 (n_4509), .B0 (n_2039), .Y(n_4309));
NAND2X1 g39917(.A (u3_mem_b2_b_34 ), .B (n_3207), .Y (n_2878));
NAND2X1 g36456(.A (n_5879), .B (n_5876), .Y (n_5877));
OAI21X1 g33775(.A0 (n_5036), .A1 (n_9105), .B0 (n_7752), .Y (n_9103));
AOI21X1 g30862(.A0 (n_12195), .A1 (n_12196), .B0 (n_11069), .Y(n_11061));
AOI21X1 g30863(.A0 (n_12064), .A1 (n_12065), .B0 (n_11059), .Y(n_11060));
NOR2X1 g30860(.A (n_10982), .B (n_11144), .Y (n_11145));
AOI21X1 g30861(.A0 (n_12193), .A1 (n_12194), .B0 (n_11069), .Y(n_11062));
AOI21X1 g30866(.A0 (n_10607), .A1 (n_10188), .B0 (n_5825), .Y(n_11056));
AOI21X1 g30867(.A0 (n_11743), .A1 (n_11744), .B0 (n_5839), .Y(n_11055));
AOI21X1 g30864(.A0 (n_10609), .A1 (n_12505), .B0 (n_11059), .Y(n_11058));
AOI21X1 g30865(.A0 (n_12793), .A1 (n_12794), .B0 (n_11059), .Y(n_11057));
NAND2X1 g39519(.A (u7_mem_b1_b_66 ), .B (n_3522), .Y (n_3124));
NAND2X1 g39518(.A (n_12369), .B (u6_mem_b0_b_108 ), .Y (n_3125));
AOI21X1 g30868(.A0 (n_12543), .A1 (n_11746), .B0 (n_5839), .Y(n_11054));
AOI21X1 g30869(.A0 (n_11749), .A1 (n_11750), .B0 (n_5839), .Y(n_11053));
NOR2X1 g35818(.A (n_740), .B (n_6752), .Y (n_6749));
NOR2X1 g35819(.A (n_495), .B (n_6752), .Y (n_6751));
MX2X1 g34141(.A (u8_mem_b0_b_111 ), .B (n_3831), .S0 (n_7490), .Y(n_8705));
MX2X1 g34140(.A (u8_mem_b0_b_110 ), .B (n_3830), .S0 (n_7490), .Y(n_8707));
MX2X1 g34143(.A (u8_mem_b0_b_113 ), .B (n_3836), .S0 (n_7490), .Y(n_8703));
MX2X1 g34142(.A (u8_mem_b0_b_112 ), .B (n_3833), .S0 (n_7490), .Y(n_8704));
MX2X1 g34145(.A (u8_mem_b0_b_114 ), .B (n_3838), .S0 (n_7490), .Y(n_8699));
MX2X1 g34144(.A (u3_mem_b0_b_113 ), .B (n_3592), .S0 (n_8700), .Y(n_8701));
MX2X1 g34147(.A (u3_mem_b0_b_114 ), .B (n_3627), .S0 (n_8700), .Y(n_8696));
MX2X1 g34146(.A (u8_mem_b0_b_115 ), .B (n_3590), .S0 (n_7490), .Y(n_8698));
MX2X1 g34148(.A (u8_mem_b0_b_116 ), .B (n_3589), .S0 (n_7490), .Y(n_9379));
INVX1 g42308(.A (u11_mem_b1_b_125 ), .Y (n_6548));
OAI21X1 g33593(.A0 (n_5078), .A1 (n_9336), .B0 (n_7960), .Y (n_9330));
INVX1 g42563(.A (n_782), .Y (n_762));
OAI21X1 g33889(.A0 (n_4881), .A1 (n_8961), .B0 (n_7635), .Y (n_8962));
OAI21X1 g33888(.A0 (n_4898), .A1 (n_8961), .B0 (n_7636), .Y (n_8963));
OAI21X1 g33885(.A0 (n_4883), .A1 (n_9038), .B0 (n_7639), .Y (n_8967));
OAI21X1 g33884(.A0 (n_5159), .A1 (n_9038), .B0 (n_7640), .Y (n_8968));
OAI21X1 g33887(.A0 (n_4882), .A1 (n_9038), .B0 (n_7637), .Y (n_8964));
OAI21X1 g33886(.A0 (n_5073), .A1 (n_9038), .B0 (n_7638), .Y (n_8965));
OAI21X1 g33881(.A0 (n_4952), .A1 (n_8971), .B0 (n_7643), .Y (n_8972));
OAI21X1 g33880(.A0 (n_5076), .A1 (n_8971), .B0 (n_7644), .Y (n_8973));
OAI21X1 g33883(.A0 (n_4884), .A1 (n_8971), .B0 (n_7641), .Y (n_8969));
OAI21X1 g33882(.A0 (n_5057), .A1 (n_8971), .B0 (n_7642), .Y (n_8970));
AOI21X1 g38020(.A0 (u7_mem_b2_b_55 ), .A1 (n_4509), .B0 (n_1948), .Y(n_4529));
NOR2X1 g40108(.A (n_2120), .B (n_2829), .Y (n_2127));
AOI21X1 g38021(.A0 (u3_mem_b2_b_43 ), .A1 (n_4533), .B0 (n_2079), .Y(n_4528));
NOR2X1 g40104(.A (n_2083), .B (n_2782), .Y (n_2130));
NAND3X1 g39111(.A (u7_mem_b0_b_92 ), .B (n_907), .C (n_1921), .Y(n_1499));
AOI21X1 g38083(.A0 (u8_mem_b2_b_33 ), .A1 (n_4491), .B0 (n_1805), .Y(n_4489));
INVX2 g32937(.A (n_9905), .Y (n_10839));
CLKBUFX3 g32934(.A (n_9818), .Y (n_10391));
BUFX3 g32933(.A (n_9674), .Y (n_9721));
NOR2X1 g40230(.A (n_2020), .B (n_2804), .Y (n_2021));
NOR2X1 g40231(.A (n_2775), .B (n_2702), .Y (n_2704));
AOI21X1 g38084(.A0 (u8_mem_b3_b_143 ), .A1 (n_3879), .B0 (n_1479), .Y(n_3878));
NOR2X1 g40233(.A (n_2713), .B (n_2829), .Y (n_2701));
AOI21X1 g38305(.A0 (u5_mem_b2_b_38 ), .A1 (n_4378), .B0 (n_1935), .Y(n_4377));
NOR2X1 g40236(.A (n_2713), .B (n_2755), .Y (n_2699));
NOR2X1 g40237(.A (n_2477), .B (n_2707), .Y (n_1827));
NOR2X1 g40238(.A (n_2775), .B (n_2716), .Y (n_2698));
NOR2X1 g40239(.A (n_2707), .B (n_1985), .Y (n_2018));
NAND2X1 g39230(.A (in_slt_399), .B (n_3415), .Y (n_3351));
NOR2X1 g39231(.A (n_5059), .B (n_2702), .Y (n_3350));
INVX1 g42560(.A (n_762), .Y (n_888));
AOI21X1 g38085(.A0 (u6_mem_b2_b_41 ), .A1 (n_4504), .B0 (n_1952), .Y(n_4488));
NAND2X1 g39233(.A (in_slt_404), .B (n_3415), .Y (n_3347));
NAND2X1 g32688(.A (n_265), .B (n_10645), .Y (n_11963));
NAND2X1 g32689(.A (n_375), .B (n_10645), .Y (n_11977));
NOR2X1 g40355(.A (n_2761), .B (n_2772), .Y (n_2657));
NOR2X1 g40354(.A (n_2470), .B (n_2735), .Y (n_1943));
NOR2X1 g40353(.A (n_2775), .B (n_2792), .Y (n_2658));
MX2X1 g35971(.A (n_461), .B (n_6510), .S0 (n_5409), .Y (n_6670));
MX2X1 g38658(.A (u5_mem_b0_b_112 ), .B (wb_din_682), .S0 (n_3720), .Y(n_3717));
NOR2X1 g39137(.A (n_2782), .B (n_1488), .Y (n_1495));
NAND2X1 g32680(.A (n_201), .B (n_10645), .Y (n_11959));
NAND2X1 g32681(.A (n_217), .B (n_10645), .Y (n_11997));
NAND2X1 g32682(.A (n_363), .B (n_10645), .Y (n_11961));
NAND2X1 g39237(.A (n_1404), .B (u3_rp_b3_b ), .Y (n_4836));
INVX2 g32685(.A (n_9642), .Y (n_9777));
NOR2X1 g40359(.A (n_2775), .B (n_2720), .Y (n_2653));
OR2X1 g32687(.A (n_1203), .B (n_9514), .Y (n_9642));
AOI21X1 g38062(.A0 (u8_mem_b2_b_45 ), .A1 (n_4499), .B0 (n_2004), .Y(n_4500));
AOI21X1 g38063(.A0 (u6_mem_b2_b_43 ), .A1 (n_4504), .B0 (n_1984), .Y(n_4498));
AOI21X1 g38060(.A0 (u7_mem_b2_b_48 ), .A1 (n_4509), .B0 (n_1964), .Y(n_4501));
AOI21X1 g38066(.A0 (u8_mem_b3_b_136 ), .A1 (n_3879), .B0 (n_1423), .Y(n_3884));
AOI21X1 g38064(.A0 (u7_mem_b1_b_77 ), .A1 (n_5118), .B0 (n_2722), .Y(n_5128));
AOI21X1 g38065(.A0 (u3_mem_b3_b_123 ), .A1 (n_5133), .B0 (n_3067), .Y(n_5127));
AOI21X1 g38068(.A0 (u7_mem_b2_b_29 ), .A1 (n_4540), .B0 (n_2001), .Y(n_4496));
AOI21X1 g38069(.A0 (u3_mem_b3_b_130 ), .A1 (n_5133), .B0 (n_3512), .Y(n_5126));
NAND2X1 g37467(.A (u13_ints_r_b15_b ), .B (n_3985), .Y (n_2578));
AOI21X1 g38224(.A0 (u4_mem_b3_b_125 ), .A1 (n_5106), .B0 (n_2953), .Y(n_5072));
INVX1 g42441(.A (u9_mem_b1_b_148 ), .Y (n_2506));
MX2X1 g38686(.A (u6_mem_b0_b_108 ), .B (wb_din_678), .S0 (n_3632), .Y(n_3674));
MX2X1 g38687(.A (u6_mem_b0_b_113 ), .B (wb_din_683), .S0 (n_3632), .Y(n_3671));
MX2X1 g38684(.A (u6_mem_b0_b_105 ), .B (wb_din_675), .S0 (n_3632), .Y(n_3676));
MX2X1 g38685(.A (u6_mem_b0_b_106 ), .B (wb_din_676), .S0 (n_3632), .Y(n_3675));
MX2X1 g38682(.A (u6_mem_b0_b_103 ), .B (wb_din_673), .S0 (n_3632), .Y(n_3679));
MX2X1 g38683(.A (u7_mem_b0_b_100 ), .B (wb_din_670), .S0 (n_3622), .Y(n_3677));
MX2X1 g38680(.A (u6_mem_b0_b_100 ), .B (wb_din_670), .S0 (n_813), .Y(n_3682));
MX2X1 g38681(.A (u6_mem_b0_b_102 ), .B (wb_din_672), .S0 (n_3632), .Y(n_3681));
MX2X1 g38688(.A (u6_mem_b0_b_116 ), .B (wb_din_686), .S0 (n_3632), .Y(n_3670));
INVX2 g41332(.A (n_851), .Y (n_1060));
INVX8 g41334(.A (n_1060), .Y (n_3826));
AND2X1 g41339(.A (n_58), .B (n_178), .Y (n_851));
NAND2X1 g36303(.A (n_2624), .B (n_2621), .Y (n_2625));
NAND2X1 g36305(.A (n_4081), .B (n_2617), .Y (n_4087));
NAND2X1 g36304(.A (n_1291), .B (n_1290), .Y (n_1292));
NAND2X1 g36307(.A (n_6821), .B (n_12626), .Y (n_5941));
NAND2X1 g36309(.A (n_6266), .B (n_6824), .Y (n_6326));
NAND2X1 g40825(.A (n_5588), .B (n_802), .Y (n_8205));
NAND2X1 g40824(.A (n_544), .B (oc2_cfg_986), .Y (n_806));
NOR2X1 g40827(.A (n_145), .B (u4_rp_b3_b ), .Y (n_712));
NOR2X1 g40826(.A (n_12634), .B (u7_rp_b3_b ), .Y (n_650));
MX2X1 g31308(.A (n_5666), .B (n_1615), .S0 (n_9721), .Y (n_10440));
AOI21X1 g31658(.A0 (n_7164), .A1 (n_1130), .B0 (n_9501), .Y (n_9502));
AOI21X1 g31659(.A0 (n_7163), .A1 (n_1116), .B0 (n_9499), .Y (n_9500));
MX2X1 g31304(.A (n_5664), .B (n_1628), .S0 (n_10537), .Y (n_10444));
MX2X1 g31305(.A (n_5655), .B (n_1755), .S0 (n_10537), .Y (n_10443));
AOI21X1 g31654(.A0 (n_7166), .A1 (n_1122), .B0 (n_12847), .Y(n_9506));
AOI21X1 g31655(.A0 (n_7289), .A1 (n_1127), .B0 (n_12845), .Y(n_9563));
NAND2X1 g31653(.A (n_1700), .B (n_10054), .Y (n_9994));
NAND2X1 g31650(.A (n_10985), .B (n_5772), .Y (n_9842));
OR2X1 g31651(.A (n_10327), .B (n_771), .Y (n_9996));
INVX1 g41484(.A (n_12801), .Y (n_1071));
BUFX3 g41486(.A (n_1072), .Y (n_5656));
NOR2X1 g41480(.A (u13_ints_r_b12_b ), .B (n_676), .Y (n_677));
NOR2X1 g41481(.A (u13_ints_r_b3_b ), .B (n_616), .Y (n_617));
INVX1 g41483(.A (n_1071), .Y (n_1384));
INVX1 g42220(.A (u11_mem_b0_b_175 ), .Y (n_1605));
OAI21X1 g45530(.A0 (n_6079), .A1 (n_11934), .B0 (n_12532), .Y(n_12136));
INVX1 g42566(.A (u9_mem_b0_b_174 ), .Y (n_1701));
INVX1 g42683(.A (u9_mem_b1_b_138 ), .Y (n_356));
INVX1 g42682(.A (u10_mem_b2_b_95 ), .Y (n_6021));
INVX1 g42681(.A (u11_mem_b1_b_148 ), .Y (n_1584));
INVX1 g42680(.A (n_8197), .Y (n_598));
NOR2X1 g40351(.A (n_832), .B (n_931), .Y (n_1199));
AOI21X1 g40350(.A0 (ic2_cfg_1044), .A1 (n_209), .B0(u14_u8_full_empty_r), .Y (n_811));
INVX1 g42466(.A (dma_req_o_b3_b), .Y (n_118));
INVX1 g42465(.A (crac_wr), .Y (n_324));
INVX1 g42464(.A (n_8550), .Y (n_465));
INVX1 g42461(.A (u9_rp_b1_b ), .Y (n_53));
XOR2X1 g35487(.A (u9_wp_b3_b ), .B (n_1557), .Y (n_4845));
NAND4X1 g35485(.A (n_5249), .B (wb_cyc_i), .C (n_303), .D (wb_stb_i),.Y (n_6051));
INVX1 g35484(.A (n_6051), .Y (n_6716));
MX2X1 g35483(.A (n_1818), .B (u2_res_cnt_b2_b ), .S0 (n_5632), .Y(n_4846));
AOI21X1 g35482(.A0 (u10_rp_b2_b ), .A1 (i4_re), .B0 (n_6711), .Y(n_7145));
AOI21X1 g35481(.A0 (u11_rp_b2_b ), .A1 (i6_re), .B0 (n_6715), .Y(n_7146));
NAND2X1 g34324(.A (n_6705), .B (n_7473), .Y (n_8243));
NAND2X1 g45897(.A (n_12169), .B (u6_mem_b1_b_73 ), .Y (n_12625));
NAND2X1 g39308(.A (u3_mem_b2_b_35 ), .B (n_3207), .Y (n_3289));
NOR2X1 g34327(.A (n_1424), .B (n_8141), .Y (n_8241));
XOR2X1 g35489(.A (u10_wp_b3_b ), .B (n_1559), .Y (n_4844));
AOI21X1 g35488(.A0 (i4_dout_617), .A1 (n_7468), .B0 (n_7133), .Y(n_7329));
NAND2X1 g36930(.A (n_1665), .B (n_1664), .Y (n_4028));
NAND2X1 g34326(.A (n_6677), .B (n_7472), .Y (n_8242));
NAND2X1 g36936(.A (n_2531), .B (n_1236), .Y (n_4812));
NAND2X1 g36937(.A (n_1654), .B (n_1652), .Y (n_4024));
NAND2X1 g36934(.A (n_1660), .B (n_1658), .Y (n_4026));
NAND2X1 g36935(.A (n_1656), .B (n_1655), .Y (n_4025));
OAI21X1 g33440(.A0 (n_4532), .A1 (n_8393), .B0 (n_8138), .Y (n_8424));
OAI21X1 g33443(.A0 (n_3856), .A1 (n_8457), .B0 (n_8133), .Y (n_8420));
NAND2X1 g34322(.A (u3_mem_b3_b_127 ), .B (n_8141), .Y (n_8075));
NAND2X1 g39375(.A (u3_mem_b2_b_47 ), .B (n_12619), .Y (n_3227));
NAND2X1 g34329(.A (u3_mem_b2_b ), .B (n_8101), .Y (n_8071));
NAND2X1 g34328(.A (n_6676), .B (n_7461), .Y (n_8238));
NOR2X1 g39374(.A (n_3332), .B (n_2684), .Y (n_3228));
NAND2X1 g34777(.A (u7_mem_b2_b_34 ), .B (n_7651), .Y (n_7657));
NAND2X1 g34688(.A (u6_mem_b3_b_151 ), .B (n_7758), .Y (n_7736));
NAND2X1 g34689(.A (u6_mem_b3_b_152 ), .B (n_7758), .Y (n_7735));
NAND2X1 g34682(.A (u6_mem_b3_b_146 ), .B (n_7758), .Y (n_7742));
NAND2X1 g34683(.A (u6_mem_b3_b_147 ), .B (n_7758), .Y (n_7741));
NAND2X1 g34680(.A (u6_mem_b3_b_144 ), .B (n_7758), .Y (n_7744));
NAND2X1 g34681(.A (u6_mem_b3_b_145 ), .B (n_7758), .Y (n_7743));
NAND2X1 g34686(.A (u6_mem_b3_b_150 ), .B (n_7758), .Y (n_7738));
NAND2X1 g34687(.A (u6_mem_b3_b_123 ), .B (n_7758), .Y (n_7737));
NAND2X1 g34684(.A (u6_mem_b3_b_148 ), .B (n_7758), .Y (n_7740));
NAND2X1 g34685(.A (u6_mem_b3_b_149 ), .B (n_7758), .Y (n_7739));
AOI21X1 g38247(.A0 (u6_mem_b3_b_148 ), .A1 (n_5059), .B0 (n_3220), .Y(n_5060));
NAND2X1 g39376(.A (u7_mem_b1_b_86 ), .B (n_4130), .Y (n_4198));
OAI21X1 g33434(.A0 (n_3885), .A1 (n_8433), .B0 (n_8146), .Y (n_8431));
OAI21X1 g33435(.A0 (n_4348), .A1 (n_8101), .B0 (n_8144), .Y (n_8430));
OAI21X1 g33436(.A0 (n_3854), .A1 (n_8930), .B0 (n_8143), .Y (n_8428));
OAI21X1 g33437(.A0 (n_4534), .A1 (n_8440), .B0 (n_8142), .Y (n_8427));
NAND2X1 g34350(.A (u4_mem_b1_b_70 ), .B (n_7984), .Y (n_8054));
NAND2X1 g34351(.A (n_6688), .B (n_7467), .Y (n_8233));
OAI21X1 g33432(.A0 (n_3883), .A1 (n_8433), .B0 (n_8148), .Y (n_8434));
OAI21X1 g33433(.A0 (n_4537), .A1 (n_8101), .B0 (n_8071), .Y (n_8432));
NAND2X1 g38829(.A (u6_mem_b3_b_145 ), .B (n_2465), .Y (n_2448));
NAND2X1 g34358(.A (u4_mem_b1_b_76 ), .B (n_7984), .Y (n_8045));
NAND2X1 g34359(.A (u4_mem_b1_b_77 ), .B (n_7984), .Y (n_8044));
NAND2X1 g34428(.A (u4_mem_b2_b_36 ), .B (n_7984), .Y (n_7988));
NAND2X1 g34429(.A (u4_mem_b2_b_37 ), .B (n_7984), .Y (n_7987));
INVX1 g42323(.A (u9_mem_b3_b_81 ), .Y (n_5302));
NAND2X1 g39371(.A (n_12679), .B (u5_mem_b0_b_116 ), .Y (n_3231));
AOI21X1 g38479(.A0 (u7_mem_b1_b_75 ), .A1 (n_5069), .B0 (n_2674), .Y(n_4901));
AOI21X1 g38478(.A0 (u7_mem_b1_b ), .A1 (n_5069), .B0 (n_2671), .Y(n_4902));
AOI21X1 g38475(.A0 (u8_mem_b3_b_137 ), .A1 (n_3879), .B0 (n_1322), .Y(n_3847));
AOI21X1 g38474(.A0 (u7_mem_b1_b_69 ), .A1 (n_5118), .B0 (n_2692), .Y(n_4905));
AOI21X1 g38477(.A0 (u7_mem_b1_b_73 ), .A1 (n_5069), .B0 (n_2699), .Y(n_4903));
AOI21X1 g38476(.A0 (u7_mem_b1_b_71 ), .A1 (n_5118), .B0 (n_2701), .Y(n_4904));
AOI21X1 g38471(.A0 (u7_mem_b3_b_132 ), .A1 (n_4961), .B0 (n_3079), .Y(n_4907));
AOI21X1 g38470(.A0 (n_1484), .A1 (n_760), .B0 (n_1485), .Y (n_3849));
AOI21X1 g38473(.A0 (u3_mem_b2_b_52 ), .A1 (n_4533), .B0 (n_2121), .Y(n_4320));
AOI21X1 g38472(.A0 (u6_mem_b1_b_68 ), .A1 (n_5112), .B0 (n_2659), .Y(n_4906));
AOI21X1 g38242(.A0 (u8_mem_b1_b_89 ), .A1 (n_4387), .B0 (n_2005), .Y(n_4393));
INVX4 g40686(.A (n_1180), .Y (n_2067));
NAND2X2 g39373(.A (n_3259), .B (u5_mem_b0_b_104 ), .Y (n_3229));
AOI21X1 g38219(.A0 (u4_mem_b3_b_151 ), .A1 (n_5106), .B0 (n_2865), .Y(n_5077));
XOR2X1 g38218(.A (n_1446), .B (n_507), .Y (n_2487));
NAND2X1 g39372(.A (u5_mem_b1_b_73 ), .B (n_3257), .Y (n_12805));
AOI21X1 g38211(.A0 (u4_mem_b3_b_147 ), .A1 (n_5102), .B0 (n_2928), .Y(n_5084));
AOI21X1 g38210(.A0 (u8_mem_b1_b_84 ), .A1 (n_4502), .B0 (n_2156), .Y(n_4400));
AOI21X1 g38213(.A0 (u4_mem_b3_b_148 ), .A1 (n_5106), .B0 (n_3246), .Y(n_5082));
AOI21X1 g38212(.A0 (u7_mem_b1_b_60 ), .A1 (n_5069), .B0 (n_2673), .Y(n_5083));
AOI21X1 g38214(.A0 (u4_mem_b3_b_149 ), .A1 (n_5106), .B0 (n_2958), .Y(n_5081));
AOI21X1 g38217(.A0 (u4_mem_b3_b_123 ), .A1 (n_5102), .B0 (n_2877), .Y(n_5078));
INVX1 g42637(.A (u10_mem_b2_b_98 ), .Y (n_6668));
NAND2X1 g45545(.A (n_6769), .B (u7_rp_b0_b ), .Y (n_12152));
AOI21X1 g32744(.A0 (n_6160), .A1 (n_5804), .B0 (n_9873), .Y(n_10574));
INVX4 g32747(.A (n_9685), .Y (n_9860));
NAND2X1 g45546(.A (n_12634), .B (n_6264), .Y (n_12153));
NAND2X1 g32741(.A (n_82), .B (n_10605), .Y (n_11736));
NAND2X1 g32740(.A (n_19), .B (n_10583), .Y (n_11626));
NAND2X1 g32742(.A (n_383), .B (n_10583), .Y (n_11630));
INVX1 g42635(.A (u10_mem_b3_b_75 ), .Y (n_5575));
OR2X1 g32749(.A (n_9641), .B (n_9564), .Y (n_9685));
CLKBUFX3 g45914(.A (n_12662), .Y (n_12645));
NAND2X1 g37867(.A (n_4120), .B (n_2970), .Y (n_5202));
NAND2X1 g45447(.A (n_12026), .B (n_12027), .Y (n_11855));
CLKBUFX3 g45912(.A (n_12662), .Y (n_12641));
AOI22X1 g37864(.A0 (n_2502), .A1 (n_6400), .B0 (n_6540), .B1(n_1859), .Y (n_1568));
NOR2X1 g39281(.A (n_4961), .B (n_2684), .Y (n_3324));
AOI22X1 g45448(.A0 (u7_mem_b2_b_34 ), .A1 (n_12641), .B0 (n_2330), .B1(u7_mem_b0_b_96 ), .Y (n_12027));
INVX1 g42565(.A (u6_rp_b2_b ), .Y (n_192));
AOI22X1 g45449(.A0 (u7_mem_b3_b_127 ), .A1 (n_1538), .B0 (n_11853),.B1 (u7_mem_b1_b_65 ), .Y (n_12026));
NOR2X1 g40857(.A (n_8197), .B (n_804), .Y (n_9695));
NAND2X1 g36442(.A (n_11925), .B (n_12531), .Y (n_6793));
MX2X1 g36115(.A (n_6442), .B (n_6441), .S0 (n_6649), .Y (n_6443));
MX2X1 g36116(.A (n_6439), .B (n_6442), .S0 (n_5409), .Y (n_6440));
NAND2X1 g36441(.A (n_6794), .B (u4_rp_b0_b ), .Y (n_11542));
MX2X1 g36110(.A (n_501), .B (n_6011), .S0 (n_6475), .Y (n_5973));
MX2X1 g36111(.A (n_509), .B (n_6925), .S0 (n_6898), .Y (n_6871));
MX2X1 g36112(.A (n_406), .B (n_6008), .S0 (n_6475), .Y (n_5971));
MX2X1 g36113(.A (n_6448), .B (n_6497), .S0 (n_932), .Y (n_6449));
NAND2X1 g39037(.A (in_slt_404), .B (n_2368), .Y (n_4778));
NAND2X1 g36448(.A (n_6244), .B (n_6259), .Y (n_6245));
MX2X1 g36118(.A (n_6434), .B (n_6486), .S0 (n_5312), .Y (n_6435));
MX2X1 g36119(.A (n_6431), .B (n_6483), .S0 (n_5312), .Y (n_6432));
NAND2X1 g39592(.A (u6_mem_b2_b_41 ), .B (n_2285), .Y (n_2278));
AND2X1 g41504(.A (n_564), .B (n_802), .Y (n_8207));
AOI21X1 g35573(.A0 (n_6825), .A1 (n_6123), .B0 (n_7324), .Y (n_7327));
INVX1 g41501(.A (n_1127), .Y (n_1381));
NOR2X1 g35571(.A (i3_re), .B (u9_rp_b0_b ), .Y (n_6714));
NAND3X1 g30050(.A (n_9769), .B (n_9601), .C (n_9661), .Y (n_10092));
OR2X1 g41503(.A (n_510), .B (n_458), .Y (n_854));
NAND2X1 g39014(.A (n_12389), .B (u4_mem_b0_b_116 ), .Y (n_3516));
INVX1 g41502(.A (n_854), .Y (n_1127));
OAI21X1 g30056(.A0 (n_9563), .A1 (n_9647), .B0 (n_9838), .Y(n_10401));
OAI21X1 g30055(.A0 (n_9506), .A1 (n_9591), .B0 (n_9756), .Y(n_10090));
AOI21X1 g35574(.A0 (n_6834), .A1 (n_6127), .B0 (n_7324), .Y (n_7326));
INVX4 g45894(.A (n_12620), .Y (n_12621));
INVX1 g41800(.A (n_593), .Y (n_5225));
INVX2 g41801(.A (wb_addr_i_b5_b), .Y (n_593));
NAND2X1 g39469(.A (n_12825), .B (u3_mem_b0_b_113 ), .Y (n_3159));
OAI21X1 g30059(.A0 (n_9502), .A1 (n_9587), .B0 (n_9754), .Y(n_10088));
NAND2X1 g39468(.A (u5_mem_b2_b_48 ), .B (n_12823), .Y (n_1791));
AOI21X1 g35578(.A0 (n_5586), .A1 (n_3976), .B0 (n_7353), .Y (n_7133));
AND2X1 g41723(.A (n_706), .B (n_751), .Y (n_813));
INVX1 g41804(.A (u9_mem_b0_b_175 ), .Y (n_1704));
MX2X1 g31130(.A (n_6903), .B (n_6902), .S0 (n_10235), .Y (n_10269));
NAND2X1 g39465(.A (u7_mem_b1_b_77 ), .B (n_3522), .Y (n_3161));
NAND2X1 g39464(.A (n_12369), .B (u6_mem_b0_b_112 ), .Y (n_3162));
INVX1 g41807(.A (u9_mem_b0_b_166 ), .Y (n_6864));
NAND2X1 g39467(.A (n_11789), .B (u8_mem_b0_b_114 ), .Y (n_3160));
INVX1 g42097(.A (u9_mem_b0_b_179 ), .Y (n_2507));
NAND2X1 g39466(.A (u4_mem_b2_b ), .B (n_12079), .Y (n_1786));
INVX1 g42090(.A (n_8188), .Y (n_670));
INVX1 g42091(.A (u10_mem_b2_b_107 ), .Y (n_98));
NAND2X1 g39461(.A (u4_mem_b1_b_71 ), .B (n_12250), .Y (n_11657));
INVX1 g42098(.A (u10_mem_b0_b_163 ), .Y (n_6375));
NOR2X1 g39460(.A (n_3332), .B (n_2707), .Y (n_3164));
AOI21X1 g38026(.A0 (u3_mem_b1_b_71 ), .A1 (n_5148), .B0 (n_2830), .Y(n_5144));
NAND2X1 g39463(.A (u5_mem_b2_b_49 ), .B (n_12823), .Y (n_2297));
NOR2X1 g39462(.A (n_3453), .B (n_2735), .Y (n_3163));
AOI21X1 g38024(.A0 (u8_mem_b1_b_90 ), .A1 (n_4502), .B0 (n_2351), .Y(n_4527));
AOI21X1 g38022(.A0 (u7_mem_b3_b_129 ), .A1 (n_5145), .B0 (n_3065), .Y(n_5146));
AND2X1 g41673(.A (n_746), .B (n_705), .Y (n_913));
INVX2 g41672(.A (n_913), .Y (n_1108));
NAND2X1 g39539(.A (u7_mem_b1_b_68 ), .B (n_3522), .Y (n_3105));
NAND2X1 g39538(.A (u7_mem_b2_b_33 ), .B (n_12654), .Y (n_3106));
NAND3X1 g30848(.A (n_8848), .B (n_1887), .C (n_7533), .Y (n_9490));
AOI21X1 g30849(.A0 (n_10623), .A1 (n_10206), .B0 (n_11144), .Y(n_11073));
INVX1 g41674(.A (n_12144), .Y (n_7324));
AOI21X1 g30844(.A0 (n_11962), .A1 (n_11963), .B0 (n_5827), .Y(n_11077));
AOI21X1 g30845(.A0 (n_11976), .A1 (n_11977), .B0 (n_11086), .Y(n_11076));
AOI21X1 g30846(.A0 (n_10626), .A1 (n_10209), .B0 (n_11069), .Y(n_11075));
AOI21X1 g30840(.A0 (n_11956), .A1 (n_11957), .B0 (n_11083), .Y(n_11081));
AOI21X1 g30841(.A0 (n_11958), .A1 (n_11959), .B0 (n_11083), .Y(n_11080));
AOI21X1 g30842(.A0 (n_11996), .A1 (n_11997), .B0 (n_11083), .Y(n_11079));
AOI21X1 g30843(.A0 (n_11960), .A1 (n_11961), .B0 (n_11083), .Y(n_11078));
AOI21X1 g38246(.A0 (u8_mem_b2_b_51 ), .A1 (n_4499), .B0 (n_2062), .Y(n_4390));
MX2X1 g34169(.A (u3_mem_b0_b_95 ), .B (n_3771), .S0 (n_8700), .Y(n_9368));
MX2X1 g34168(.A (u3_mem_b0_b_94 ), .B (n_3575), .S0 (n_8700), .Y(n_8682));
INVX1 g42324(.A (u10_mem_b1_b_139 ), .Y (n_249));
INVX1 g42325(.A (u11_mem_b1_b_142 ), .Y (n_1614));
MX2X1 g37215(.A (u10_mem_b2_b_112 ), .B (n_5355), .S0 (n_5341), .Y(n_5377));
MX2X1 g34163(.A (u8_mem_b0_b_98 ), .B (n_3649), .S0 (n_7490), .Y(n_8687));
MX2X1 g34162(.A (u8_mem_b0_b_97 ), .B (n_3570), .S0 (n_7490), .Y(n_8688));
MX2X1 g34161(.A (u8_mem_b0_b_96 ), .B (n_3750), .S0 (n_7490), .Y(n_8689));
MX2X1 g34160(.A (u3_mem_b0_b_119 ), .B (n_3582), .S0 (n_8700), .Y(n_9369));
MX2X1 g34167(.A (u3_mem_b0_b_93 ), .B (n_3744), .S0 (n_7423), .Y(n_8684));
MX2X1 g34166(.A (u3_mem_b0_b_121 ), .B (n_3577), .S0 (n_7423), .Y(n_8250));
MX2X1 g34165(.A (u3_mem_b0_b_120 ), .B (n_3579), .S0 (n_8700), .Y(n_8685));
MX2X1 g34164(.A (u8_mem_b0_b_99 ), .B (n_3580), .S0 (n_7490), .Y(n_8686));
AOI21X1 g38245(.A0 (u8_mem_b1_b_73 ), .A1 (n_4502), .B0 (n_1988), .Y(n_4391));
NAND2X1 g37746(.A (n_3240), .B (n_3238), .Y (n_4596));
AOI21X1 g38243(.A0 (u3_mem_b2_b_58 ), .A1 (n_4519), .B0 (n_2086), .Y(n_4392));
NAND2X1 g39797(.A (n_3252), .B (u7_mem_b0_b_118 ), .Y (n_2952));
NOR2X1 g39796(.A (n_3486), .B (n_2794), .Y (n_2953));
NOR2X1 g39794(.A (n_3089), .B (n_2792), .Y (n_2954));
NAND2X1 g39793(.A (u6_mem_b2_b_52 ), .B (n_3423), .Y (n_2955));
NAND2X1 g37744(.A (n_3176), .B (n_3071), .Y (n_4597));
NAND2X1 g39791(.A (n_2330), .B (u7_mem_b0_b_105 ), .Y (n_2331));
NAND2X1 g39790(.A (u7_mem_b1_b_74 ), .B (n_4130), .Y (n_4125));
MX2X1 g37213(.A (u10_mem_b2_b_109 ), .B (n_5290), .S0 (n_5424), .Y(n_5379));
NOR2X1 g39799(.A (n_3486), .B (n_2792), .Y (n_2951));
NAND2X1 g39798(.A (n_2491), .B (u7_mem_b0_b_106 ), .Y (n_2200));
NOR2X1 g36612(.A (n_2610), .B (n_2587), .Y (n_4828));
NAND2X1 g36611(.A (n_5709), .B (n_6091), .Y (n_6140));
NAND2X1 g36610(.A (n_6142), .B (n_6141), .Y (n_6143));
OAI21X1 g36616(.A0 (n_4629), .A1 (n_5200), .B0 (n_784), .Y (n_6139));
OR2X1 g36343(.A (n_1290), .B (n_4633), .Y (n_2619));
INVX2 g40781(.A (n_945), .Y (n_1172));
NAND2X2 g40782(.A (n_627), .B (u3_wp_b1_b ), .Y (n_945));
BUFX3 g40783(.A (n_937), .Y (n_4499));
INVX8 g40786(.A (n_1129), .Y (n_1985));
INVX1 g40787(.A (n_1129), .Y (n_2137));
NAND2X1 g45709(.A (n_12641), .B (u7_mem_b2_b_47 ), .Y (n_12410));
NAND2X1 g31641(.A (n_5357), .B (n_10010), .Y (n_10003));
NAND2X1 g39868(.A (u3_mem_b1_b_85 ), .B (n_3316), .Y (n_2911));
NAND2X1 g45457(.A (dma_req_o_b8_b), .B (n_11903), .Y (n_11905));
NOR2X1 g40225(.A (n_2025), .B (n_2748), .Y (n_2026));
INVX8 g32919(.A (n_9820), .Y (n_10513));
INVX1 g45456(.A (dma_ack_i_b8_b), .Y (n_11903));
NOR2X1 g40258(.A (n_2735), .B (n_2137), .Y (n_2004));
NOR2X1 g40259(.A (n_945), .B (n_2684), .Y (n_2003));
NOR2X1 g40252(.A (n_2096), .B (n_2691), .Y (n_2010));
NOR2X1 g40253(.A (n_867), .B (n_2772), .Y (n_2476));
NOR2X1 g40250(.A (n_2099), .B (n_2767), .Y (n_2012));
NOR2X1 g40251(.A (n_2041), .B (n_2702), .Y (n_2011));
NOR2X1 g40256(.A (n_2006), .B (n_2716), .Y (n_2007));
NOR2X1 g40257(.A (n_2864), .B (n_2057), .Y (n_2005));
NOR2X1 g40254(.A (n_2702), .B (n_2008), .Y (n_2009));
NOR2X1 g40255(.A (n_2721), .B (n_2818), .Y (n_2693));
NAND2X1 g45455(.A (u16_u8_dma_req_r1), .B (n_11903), .Y (n_11904));
CLKBUFX3 g45974(.A (n_12743), .Y (n_12744));
INVX2 g45975(.A (n_12742), .Y (n_12743));
NAND2X1 g45976(.A (n_521), .B (u4_rp_b2_b ), .Y (n_12742));
INVX1 g45977(.A (n_12743), .Y (n_12747));
INVX2 g45970(.A (n_602), .Y (n_12738));
NAND4X1 g45971(.A (n_12739), .B (n_12740), .C (n_12741), .D(n_12745), .Y (n_12746));
NAND2X1 g45972(.A (n_12389), .B (u4_mem_b0_b_103 ), .Y (n_12739));
NAND2X1 g45973(.A (n_12744), .B (u4_mem_b3_b_134 ), .Y (n_12745));
NAND4X1 g45978(.A (n_12748), .B (n_12749), .C (n_12750), .D(n_12754), .Y (n_12755));
NAND2X1 g45979(.A (n_12825), .B (u3_mem_b0_b_104 ), .Y (n_12748));
OR2X1 g40331(.A (n_910), .B (n_1484), .Y (n_1449));
NOR2X1 g40330(.A (n_2775), .B (n_2782), .Y (n_2662));
NOR2X1 g40333(.A (n_2773), .B (n_2707), .Y (n_2661));
NOR2X1 g40332(.A (n_2189), .B (n_2831), .Y (n_1959));
NOR2X1 g40335(.A (n_821), .B (n_2772), .Y (n_1958));
NOR2X1 g40334(.A (n_2761), .B (n_2729), .Y (n_2660));
NOR2X1 g40337(.A (n_2732), .B (n_2008), .Y (n_1956));
NOR2X1 g40336(.A (n_2470), .B (n_2741), .Y (n_1957));
NOR2X1 g40339(.A (n_2133), .B (n_2729), .Y (n_1954));
NOR2X1 g40338(.A (n_2083), .B (n_2763), .Y (n_1955));
AOI21X1 g38048(.A0 (u4_mem_b1_b_87 ), .A1 (n_4507), .B0 (n_2146), .Y(n_4508));
AOI21X1 g38049(.A0 (u3_mem_b3_b_134 ), .A1 (n_5138), .B0 (n_2985), .Y(n_5139));
AOI21X1 g38044(.A0 (u3_mem_b2_b_35 ), .A1 (n_4519), .B0 (n_1941), .Y(n_4512));
AOI21X1 g38045(.A0 (u3_mem_b2_b_37 ), .A1 (n_4519), .B0 (n_2027), .Y(n_4511));
AOI21X1 g38046(.A0 (u8_mem_b3_b_148 ), .A1 (n_3879), .B0 (n_1476), .Y(n_3885));
AOI21X1 g38047(.A0 (u7_mem_b2_b_49 ), .A1 (n_4509), .B0 (n_1945), .Y(n_4510));
AOI21X1 g38040(.A0 (u6_mem_b2_b_46 ), .A1 (n_4544), .B0 (n_2234), .Y(n_4515));
AOI21X1 g38041(.A0 (u4_mem_b1_b_88 ), .A1 (n_4507), .B0 (n_1999), .Y(n_4514));
AOI21X1 g38042(.A0 (u6_mem_b1_b_89 ), .A1 (n_5112), .B0 (n_2762), .Y(n_5140));
AOI21X1 g38043(.A0 (u3_mem_b2_b_34 ), .A1 (n_4519), .B0 (n_2141), .Y(n_4513));
NAND2X1 g39608(.A (n_2302), .B (in_slt_433), .Y (n_4759));
OAI21X1 g33827(.A0 (n_5005), .A1 (n_9038), .B0 (n_7696), .Y (n_9039));
NOR2X1 g39605(.A (n_3453), .B (n_2772), .Y (n_3065));
NAND2X1 g37180(.A (n_4565), .B (n_2252), .Y (n_6486));
NAND2X1 g37181(.A (n_4563), .B (n_2249), .Y (n_6547));
NAND2X1 g37182(.A (n_4561), .B (n_2248), .Y (n_6483));
NAND2X1 g37183(.A (n_3894), .B (n_3020), .Y (n_5983));
OAI21X1 g37409(.A0 (u10_mem_b0_b_179 ), .A1 (n_6341), .B0 (n_5227), .Y(n_5643));
NAND2X1 g37185(.A (n_4557), .B (n_2240), .Y (n_6573));
AOI22X1 g37638(.A0 (n_365), .A1 (n_1835), .B0 (n_5369), .B1 (n_1760),.Y (n_1730));
NAND2X1 g37187(.A (n_3928), .B (n_2305), .Y (n_6570));
NAND2X1 g37188(.A (n_4550), .B (n_2334), .Y (n_6566));
AOI22X1 g37637(.A0 (n_45), .A1 (n_1859), .B0 (n_5302), .B1 (n_1760),.Y (n_1731));
AOI22X1 g37634(.A0 (n_198), .A1 (n_1835), .B0 (n_5343), .B1 (n_1760),.Y (n_1736));
NOR2X1 g39606(.A (n_3117), .B (n_2691), .Y (n_3063));
AOI22X1 g37633(.A0 (n_2502), .A1 (n_1738), .B0 (n_1737), .B1(n_1859), .Y (n_1739));
AOI22X1 g37630(.A0 (n_356), .A1 (n_1859), .B0 (n_1744), .B1 (n_1835),.Y (n_1745));
AOI22X1 g37631(.A0 (n_2502), .A1 (n_1742), .B0 (n_5294), .B1(n_1760), .Y (n_1743));
AND2X1 g41319(.A (u12_we1), .B (wb_cyc_i), .Y (n_476));
OAI21X1 g33748(.A0 (n_4525), .A1 (n_9165), .B0 (n_7780), .Y (n_9134));
OAI21X1 g33749(.A0 (n_4531), .A1 (n_9087), .B0 (n_7779), .Y (n_9133));
OAI21X1 g33746(.A0 (n_4523), .A1 (n_9087), .B0 (n_7782), .Y (n_9137));
OAI21X1 g33747(.A0 (n_4335), .A1 (n_9170), .B0 (n_7781), .Y (n_9136));
OAI21X1 g33744(.A0 (n_4505), .A1 (n_9139), .B0 (n_7784), .Y (n_9140));
OAI21X1 g33745(.A0 (n_4515), .A1 (n_9182), .B0 (n_7783), .Y (n_9138));
OAI21X1 g33742(.A0 (n_4498), .A1 (n_9165), .B0 (n_7786), .Y (n_9142));
OAI21X1 g33743(.A0 (n_4336), .A1 (n_9182), .B0 (n_7785), .Y (n_9141));
OAI21X1 g33740(.A0 (n_4488), .A1 (n_9170), .B0 (n_7788), .Y (n_9144));
OAI21X1 g33741(.A0 (n_4337), .A1 (n_9182), .B0 (n_7787), .Y (n_9143));
NAND2X1 g36329(.A (n_6239), .B (n_6318), .Y (n_6315));
NAND2X1 g36328(.A (n_5857), .B (n_6318), .Y (n_5937));
NAND2X1 g36323(.A (n_6821), .B (n_12171), .Y (n_6826));
NAND2X1 g36322(.A (n_6254), .B (n_6824), .Y (n_6322));
NAND2X1 g36321(.A (n_12530), .B (n_6824), .Y (n_6323));
NAND2X1 g36320(.A (n_6800), .B (n_145), .Y (n_11541));
NAND2X1 g36327(.A (n_6194), .B (n_6316), .Y (n_6317));
NAND2X1 g36326(.A (n_6142), .B (n_6318), .Y (n_6319));
NAND2X1 g36325(.A (n_5719), .B (n_6318), .Y (n_6320));
NAND2X1 g36324(.A (n_6824), .B (n_6246), .Y (n_6321));
NAND2X1 g31678(.A (n_1754), .B (n_10385), .Y (n_10386));
NAND2X1 g31679(.A (n_1619), .B (n_10391), .Y (n_10384));
NAND2X1 g40809(.A (n_8188), .B (n_921), .Y (n_9587));
AND2X1 g40808(.A (u11_wp_b1_b ), .B (n_520), .Y (n_995));
OR2X1 g31670(.A (n_9496), .B (n_9483), .Y (n_9654));
OR2X1 g31671(.A (n_9495), .B (n_9481), .Y (n_9651));
AND2X1 g31672(.A (n_5615), .B (ac97_rst_force), .Y (n_9494));
NAND2X1 g31673(.A (n_5632), .B (ac97_rst_force), .Y (n_9597));
NAND2X1 g31674(.A (n_1650), .B (n_10391), .Y (n_10390));
NAND2X1 g31675(.A (n_1644), .B (n_10391), .Y (n_10389));
NAND2X1 g31676(.A (n_1633), .B (n_10385), .Y (n_10388));
NAND2X1 g31677(.A (n_339), .B (n_10385), .Y (n_10387));
AOI21X1 g35847(.A0 (n_2613), .A1 (n_4718), .B0 (n_7353), .Y (n_7106));
NAND2X1 g37458(.A (n_5277), .B (crac_out_861), .Y (n_3973));
NAND2X1 g37459(.A (u13_ints_r_b4_b ), .B (n_3985), .Y (n_2582));
NAND2X1 g37980(.A (n_1386), .B (n_4148), .Y (n_5451));
NAND2X1 g37981(.A (n_2380), .B (n_3052), .Y (n_5165));
NAND2X1 g37982(.A (n_3191), .B (n_3030), .Y (n_5164));
NAND2X1 g37983(.A (n_3282), .B (n_3473), .Y (n_5163));
NAND2X1 g37456(.A (u13_ints_r_b2_b ), .B (n_3979), .Y (n_3975));
NAND2X1 g37985(.A (n_3107), .B (n_2903), .Y (n_5162));
AOI22X1 g37986(.A0 (u10_din_tmp_47), .A1 (n_3339), .B0 (n_3911), .B1(in_slt_426), .Y (n_4550));
NAND2X1 g37455(.A (u13_ints_r_b28_b ), .B (n_4726), .Y (n_2583));
NAND4X1 g33298(.A (n_5620), .B (n_1833), .C (n_8700), .D (n_822), .Y(n_9453));
INVX1 g33299(.A (n_12149), .Y (n_9943));
INVX2 g33291(.A (n_12688), .Y (n_10481));
AOI21X1 g35846(.A0 (n_2586), .A1 (n_4719), .B0 (n_7353), .Y (n_7110));
MX2X1 g37311(.A (u10_mem_b1_b_147 ), .B (n_5284), .S0 (n_5407), .Y(n_5285));
AND2X1 g41544(.A (n_319), .B (n_471), .Y (n_9719));
NOR2X1 g35845(.A (n_5404), .B (u2_bit_clk_e), .Y (n_6025));
MX2X1 g36048(.A (n_6893), .B (n_6906), .S0 (n_6898), .Y (n_6894));
NAND2X1 g36589(.A (n_6167), .B (n_12115), .Y (n_6168));
NAND2X1 g36588(.A (n_6155), .B (n_6259), .Y (n_6169));
NAND2X1 g36586(.A (n_5809), .B (n_6259), .Y (n_5810));
NOR2X1 g35844(.A (n_5403), .B (u2_bit_clk_e), .Y (n_5976));
NAND2X1 g36584(.A (n_6172), .B (n_12115), .Y (n_6173));
NAND2X1 g36583(.A (n_6174), .B (n_634), .Y (n_11986));
NAND2X1 g36582(.A (n_6176), .B (n_12664), .Y (n_6177));
NAND2X1 g36581(.A (n_11898), .B (n_12115), .Y (n_6179));
NAND2X1 g36580(.A (n_6180), .B (n_12531), .Y (n_6181));
NAND2X1 g39295(.A (u7_mem_b1_b_62 ), .B (n_4225), .Y (n_4204));
INVX1 g42669(.A (u11_mem_b2_b_99 ), .Y (n_6471));
INVX1 g42668(.A (u10_mem_b3_b_84 ), .Y (n_5352));
MX2X1 g36049(.A (n_6560), .B (n_6559), .S0 (n_5371), .Y (n_6561));
INVX1 g42664(.A (u11_mem_b0_b_152 ), .Y (n_6355));
INVX1 g42660(.A (u10_mem_b0_b_174 ), .Y (n_2550));
INVX1 g42663(.A (u11_mem_b2_b_101 ), .Y (n_6466));
NAND2X1 g39494(.A (u6_mem_b1_b_81 ), .B (n_4253), .Y (n_4182));
NAND2X1 g39496(.A (u3_mem_b2_b_36 ), .B (n_12619), .Y (n_3143));
NAND2X1 g39497(.A (n_12369), .B (u6_mem_b0_b_92 ), .Y (n_3142));
NOR2X1 g39490(.A (n_2792), .B (n_1488), .Y (n_1479));
NAND2X1 g39491(.A (u8_mem_b1_b_63 ), .B (n_12295), .Y (n_11464));
NAND2X1 g39493(.A (u8_mem_b2_b_59 ), .B (n_3441), .Y (n_3144));
NAND2X1 g39498(.A (n_2330), .B (u7_mem_b0_b_102 ), .Y (n_2294));
NAND2X1 g39499(.A (u6_mem_b1_b_61 ), .B (n_12169), .Y (n_11514));
OAI21X1 g30989(.A0 (n_4768), .A1 (n_10738), .B0 (n_10030), .Y(n_10714));
OAI21X1 g30988(.A0 (n_4765), .A1 (n_10019), .B0 (n_10031), .Y(n_10715));
OAI21X1 g30981(.A0 (n_4758), .A1 (n_10738), .B0 (n_10040), .Y(n_10725));
OAI21X1 g30980(.A0 (n_4777), .A1 (n_10747), .B0 (n_10041), .Y(n_10727));
OAI21X1 g30983(.A0 (n_4756), .A1 (n_10738), .B0 (n_9994), .Y(n_10722));
OAI21X1 g30982(.A0 (n_4775), .A1 (n_10747), .B0 (n_10038), .Y(n_10723));
OAI21X1 g30985(.A0 (n_4744), .A1 (n_10738), .B0 (n_10035), .Y(n_10719));
OAI21X1 g30984(.A0 (n_4774), .A1 (n_10747), .B0 (n_10037), .Y(n_10721));
OAI21X1 g30987(.A0 (n_4770), .A1 (n_10019), .B0 (n_10032), .Y(n_10717));
OAI21X1 g30986(.A0 (n_4773), .A1 (n_10747), .B0 (n_10034), .Y(n_10718));
NAND2X1 g35842(.A (n_5632), .B (u2_res_cnt_b0_b ), .Y (n_4094));
NAND2X1 g31582(.A (n_174), .B (n_10073), .Y (n_10074));
NAND2X1 g31583(.A (n_9), .B (n_10065), .Y (n_10072));
NAND2X1 g31580(.A (n_366), .B (n_10010), .Y (n_10076));
NAND2X1 g31581(.A (n_349), .B (n_10073), .Y (n_10075));
NOR2X1 g31586(.A (n_12339), .B (n_1096), .Y (n_10068));
NAND2X1 g31587(.A (n_2627), .B (n_10010), .Y (n_10067));
NAND2X1 g31584(.A (n_2549), .B (n_10010), .Y (n_10071));
NAND2X1 g31585(.A (n_379), .B (n_10010), .Y (n_10069));
NAND2X1 g31588(.A (n_2545), .B (n_10065), .Y (n_10066));
NAND2X1 g31589(.A (n_204), .B (n_10045), .Y (n_10064));
INVX2 g45365(.A (n_11579), .Y (n_11587));
CLKBUFX1 g45364(.A (n_11587), .Y (n_11586));
INVX2 g45366(.A (u6_rp_b1_b ), .Y (n_11579));
AOI21X1 g35352(.A0 (i4_dout_608), .A1 (n_7297), .B0 (n_7348), .Y(n_7460));
AOI21X1 g35351(.A0 (i4_dout_607), .A1 (n_7468), .B0 (n_7349), .Y(n_7461));
AOI21X1 g35350(.A0 (n_7468), .A1 (i4_dout_603), .B0 (n_7340), .Y(n_7462));
OR2X1 g35357(.A (n_7149), .B (ic0_int_set_719), .Y (n_7364));
AOI21X1 g35356(.A0 (i4_dout_604), .A1 (n_7468), .B0 (n_7339), .Y(n_7459));
NOR2X1 g35354(.A (i4_status), .B (i4_status_1032), .Y (n_7031));
NAND2X1 g39678(.A (u4_mem_b1_b_75 ), .B (n_12250), .Y (n_12828));
NOR2X1 g39679(.A (n_5059), .B (n_2686), .Y (n_2777));
OR2X1 g35359(.A (n_7018), .B (ic2_int_set_723), .Y (n_7280));
OR2X1 g35358(.A (n_7148), .B (ic1_int_set_721), .Y (n_7363));
NAND4X1 g36918(.A (n_11441), .B (n_3202), .C (n_11442), .D (n_2408),.Y (n_5863));
NAND2X1 g36919(.A (n_1837), .B (n_1653), .Y (n_4031));
INVX1 g36915(.A (n_5709), .Y (n_5710));
NAND4X1 g36916(.A (n_2243), .B (n_3206), .C (n_3205), .D (n_2439), .Y(n_5709));
INVX1 g36917(.A (n_5863), .Y (n_5558));
INVX1 g36910(.A (n_6241), .Y (n_5711));
NAND4X1 g36911(.A (n_11966), .B (n_3218), .C (n_11967), .D (n_2406),.Y (n_6241));
NAND4X1 g36912(.A (n_12857), .B (n_12858), .C (n_11482), .D (n_1336),.Y (n_5874));
NAND4X1 g36913(.A (n_3542), .B (n_3212), .C (n_2857), .D (n_2231), .Y(n_5559));
NAND2X1 g37696(.A (n_3551), .B (n_3297), .Y (n_4606));
MX2X1 g33984(.A (u4_mem_b0_b_102 ), .B (n_3799), .S0 (n_7499), .Y(n_8835));
MX2X1 g33985(.A (u4_mem_b0_b_103 ), .B (n_3797), .S0 (n_7499), .Y(n_9442));
MX2X1 g33986(.A (u4_mem_b0_b_104 ), .B (n_3796), .S0 (n_7499), .Y(n_9441));
MX2X1 g33987(.A (u4_mem_b0_b_105 ), .B (n_3795), .S0 (n_7499), .Y(n_8833));
MX2X1 g33980(.A (u3_mem_b0_b_101 ), .B (n_3811), .S0 (n_8700), .Y(n_9443));
MX2X1 g33981(.A (u4_mem_b0_b_100 ), .B (n_3802), .S0 (n_7499), .Y(n_8838));
MX2X1 g33982(.A (u4_mem_b0_b ), .B (n_3803), .S0 (n_7499), .Y(n_8837));
MX2X1 g33983(.A (u4_mem_b0_b_101 ), .B (n_3801), .S0 (n_7499), .Y(n_8836));
MX2X1 g33988(.A (u4_mem_b0_b_106 ), .B (n_3791), .S0 (n_7499), .Y(n_9440));
MX2X1 g33989(.A (u4_mem_b0_b_107 ), .B (n_3788), .S0 (n_7499), .Y(n_8832));
INVX4 g42955(.A (n_710), .Y (n_798));
NAND2X1 g34400(.A (u4_mem_b2_b_49 ), .B (n_7984), .Y (n_8005));
NAND2X1 g34401(.A (u4_mem_b2_b_50 ), .B (n_7984), .Y (n_8004));
NAND2X1 g34402(.A (u4_mem_b2_b_51 ), .B (n_7984), .Y (n_8003));
NAND2X1 g34403(.A (u4_mem_b2_b_52 ), .B (n_7984), .Y (n_8002));
AND2X1 g34404(.A (n_7287), .B (n_7443), .Y (n_7521));
INVX2 g34406(.A (n_7518), .Y (n_8643));
AOI22X1 g35704(.A0 (n_6686), .A1 (i6_dout_642), .B0 (i3_dout_580),.B1 (n_6700), .Y (n_6678));
NOR2X1 g39284(.A (n_3332), .B (n_2765), .Y (n_3318));
AOI22X1 g35706(.A0 (n_6686), .A1 (i6_dout_643), .B0 (i3_dout_581),.B1 (n_6700), .Y (n_6745));
MX2X1 g38678(.A (u7_mem_b0_b_104 ), .B (wb_din_674), .S0 (n_3622), .Y(n_3684));
NAND2X1 g39286(.A (n_2325), .B (in_slt_443), .Y (n_2329));
MX2X1 g33979(.A (u3_mem_b0_b_109 ), .B (n_3823), .S0 (n_8700), .Y(n_8839));
MX2X1 g33978(.A (u3_mem_b0_b_118 ), .B (n_3584), .S0 (n_8700), .Y(n_8841));
AOI21X1 g38189(.A0 (u4_mem_b3_b_134 ), .A1 (n_5102), .B0 (n_3307), .Y(n_5103));
AOI21X1 g38188(.A0 (u4_mem_b3_b_133 ), .A1 (n_5106), .B0 (n_3309), .Y(n_5104));
AOI22X1 g35702(.A0 (n_6686), .A1 (i6_dout_634), .B0 (n_6700), .B1(i3_dout_572), .Y (n_6681));
XOR2X1 g38181(.A (u10_rp_b2_b ), .B (n_638), .Y (n_1039));
AOI21X1 g38180(.A0 (u4_mem_b2_b_36 ), .A1 (n_4439), .B0 (n_1973), .Y(n_4408));
AOI21X1 g38183(.A0 (u6_mem_b1_b_64 ), .A1 (n_5112), .B0 (n_2753), .Y(n_5108));
AOI21X1 g38182(.A0 (u4_mem_b2_b_37 ), .A1 (n_4439), .B0 (n_2209), .Y(n_4407));
AOI21X1 g38187(.A0 (u6_mem_b2_b_35 ), .A1 (n_4504), .B0 (n_1673), .Y(n_4405));
AOI21X1 g38186(.A0 (u4_mem_b3_b_132 ), .A1 (n_5102), .B0 (n_3343), .Y(n_5105));
OAI21X1 g33975(.A0 (n_5160), .A1 (n_8393), .B0 (n_8068), .Y (n_8846));
INVX1 g42952(.A (u11_mem_b3_b ), .Y (n_6554));
INVX4 g41595(.A (n_707), .Y (n_5059));
NAND2X1 g34654(.A (u6_mem_b2_b_57 ), .B (n_7758), .Y (n_7771));
NAND2X1 g34657(.A (u6_mem_b2_b_59 ), .B (n_7758), .Y (n_7768));
NAND2X1 g38805(.A (u3_mem_b3_b_152 ), .B (n_2463), .Y (n_2456));
NAND2X1 g34656(.A (u6_mem_b2_b_58 ), .B (n_7758), .Y (n_7769));
AOI21X1 g38197(.A0 (u6_mem_b2_b_34 ), .A1 (n_4504), .B0 (n_2037), .Y(n_4403));
NAND2X1 g34651(.A (u6_mem_b2_b_54 ), .B (n_7758), .Y (n_7774));
INVX8 g41591(.A (n_1509), .Y (n_3332));
NAND2X1 g34650(.A (u6_mem_b2_b_53 ), .B (n_7758), .Y (n_7775));
OAI21X1 g33973(.A0 (n_4482), .A1 (n_8457), .B0 (n_7560), .Y (n_8850));
OAI21X1 g33972(.A0 (n_4479), .A1 (n_8868), .B0 (n_7561), .Y (n_8851));
NOR2X1 g39299(.A (n_3486), .B (n_2720), .Y (n_3299));
NOR2X1 g32769(.A (n_9365), .B (n_11128), .Y (n_9520));
MX2X1 g36164(.A (n_6366), .B (n_6510), .S0 (n_6359), .Y (n_6367));
INVX1 g32767(.A (n_12589), .Y (n_9908));
NAND3X1 g32766(.A (n_9672), .B (n_4679), .C (n_11772), .Y (n_9910));
OR2X1 g32765(.A (n_8482), .B (n_9359), .Y (n_9461));
OR2X1 g32764(.A (n_8483), .B (n_8679), .Y (n_9462));
OR2X1 g32763(.A (n_8484), .B (n_9352), .Y (n_9463));
OR2X1 g32762(.A (n_9507), .B (n_9475), .Y (n_9635));
OR2X1 g32761(.A (n_9508), .B (n_9476), .Y (n_9636));
OR2X1 g32760(.A (n_9509), .B (n_9477), .Y (n_9637));
AOI21X1 g38457(.A0 (u7_mem_b3_b_152 ), .A1 (n_4961), .B0 (n_3321), .Y(n_4912));
AOI21X1 g38456(.A0 (u8_mem_b3_b_125 ), .A1 (n_3879), .B0 (n_1414), .Y(n_3852));
AOI21X1 g38455(.A0 (u3_mem_b1_b_74 ), .A1 (n_5157), .B0 (n_2743), .Y(n_4913));
AOI21X1 g38454(.A0 (u6_mem_b3_b_129 ), .A1 (n_5100), .B0 (n_3035), .Y(n_4914));
AOI21X1 g38453(.A0 (u6_mem_b3_b_128 ), .A1 (n_5100), .B0 (n_2977), .Y(n_4915));
AOI21X1 g38452(.A0 (u6_mem_b3_b_127 ), .A1 (n_5059), .B0 (n_3318), .Y(n_4916));
AOI21X1 g38451(.A0 (u6_mem_b3_b_125 ), .A1 (n_5059), .B0 (n_3204), .Y(n_4917));
AOI21X1 g38450(.A0 (u7_mem_b1_b_70 ), .A1 (n_5118), .B0 (n_2752), .Y(n_4918));
AOI21X1 g38459(.A0 (u8_mem_b3_b_131 ), .A1 (n_3879), .B0 (n_1501), .Y(n_3851));
MX2X1 g36160(.A (n_6375), .B (n_6589), .S0 (n_6341), .Y (n_6376));
MX2X1 g36162(.A (n_6370), .B (n_6473), .S0 (n_6359), .Y (n_6371));
MX2X1 g31340(.A (n_6338), .B (n_6337), .S0 (n_10315), .Y (n_10123));
MX2X1 g31341(.A (n_6336), .B (n_6335), .S0 (n_10565), .Y (n_10411));
MX2X1 g31342(.A (n_6332), .B (n_6331), .S0 (n_10137), .Y (n_10122));
NAND2X1 g31697(.A (n_313), .B (n_10081), .Y (n_9988));
AOI21X1 g38233(.A0 (u6_mem_b2_b_58 ), .A1 (n_4504), .B0 (n_1990), .Y(n_4399));
AOI21X1 g38232(.A0 (u4_mem_b3_b_129 ), .A1 (n_5102), .B0 (n_2992), .Y(n_5065));
XOR2X1 g38231(.A (u10_wp_b3_b ), .B (n_1067), .Y (n_2486));
AOI21X1 g38230(.A0 (u8_mem_b3_b_124 ), .A1 (n_3879), .B0 (n_1478), .Y(n_3864));
AOI21X1 g38237(.A0 (u8_mem_b1_b_82 ), .A1 (n_4502), .B0 (n_2053), .Y(n_4397));
NAND2X1 g31694(.A (n_277), .B (n_10376), .Y (n_10367));
AOI21X1 g38235(.A0 (u6_mem_b2_b_59 ), .A1 (n_4544), .B0 (n_2145), .Y(n_4398));
NAND2X1 g38989(.A (u3_mem_b3_b_126 ), .B (n_1517), .Y (n_1507));
NAND2X1 g38988(.A (u3_mem_b3_b_149 ), .B (n_2463), .Y (n_2379));
AOI21X1 g38239(.A0 (u8_mem_b2_b_49 ), .A1 (n_4491), .B0 (n_2164), .Y(n_4396));
MX2X1 g31347(.A (u10_din_tmp_43), .B (in_slt_424), .S0 (n_9860), .Y(n_9872));
INVX8 g36469(.A (n_11119), .Y (n_6752));
INVX1 g41973(.A (u11_mem_b1_b_130 ), .Y (n_6515));
INVX1 g37089(.A (n_5813), .Y (n_5533));
NAND4X1 g37088(.A (n_11447), .B (n_11448), .C (n_2338), .D (n_2455),.Y (n_5898));
XOR2X1 g40379(.A (n_798), .B (n_1033), .Y (n_6047));
INVX4 g42718(.A (n_862), .Y (n_5839));
MX2X1 g38712(.A (u6_mem_b0_b_119 ), .B (wb_din_689), .S0 (n_3632), .Y(n_3633));
INVX1 g42291(.A (n_8536), .Y (n_175));
MX2X1 g38713(.A (u7_mem_b0_b_96 ), .B (wb_din_666), .S0 (n_3622), .Y(n_3631));
INVX1 g43011(.A (u10_mem_b1_b_125 ), .Y (n_6406));
MX2X1 g38676(.A (u5_mem_b0_b_96 ), .B (wb_din_666), .S0 (n_3720), .Y(n_3688));
NAND2X1 g34382(.A (u4_mem_b1_b_66 ), .B (n_7984), .Y (n_8021));
NAND2X1 g37845(.A (n_4182), .B (n_3162), .Y (n_12054));
AOI22X1 g37844(.A0 (n_6445), .A1 (n_1575), .B0 (n_6417), .B1(n_1831), .Y (n_1578));
AOI22X1 g37847(.A0 (n_6439), .A1 (n_1575), .B0 (n_6441), .B1(n_1831), .Y (n_1576));
AOI22X1 g37846(.A0 (n_1756), .A1 (n_6353), .B0 (n_6490), .B1(n_1643), .Y (n_1577));
AOI22X1 g37841(.A0 (n_1756), .A1 (n_1581), .B0 (n_1580), .B1(n_1643), .Y (n_1582));
AOI22X1 g37840(.A0 (n_190), .A1 (n_1575), .B0 (n_5508), .B1 (n_1831),.Y (n_1583));
AOI22X1 g37843(.A0 (u10_din_tmp1), .A1 (n_2302), .B0 (n_3911), .B1(in_slt_420), .Y (n_2521));
NAND2X1 g37849(.A (n_2466), .B (n_3094), .Y (n_12057));
AOI22X1 g37848(.A0 (n_1756), .A1 (n_6351), .B0 (n_6545), .B1(n_1643), .Y (n_1574));
MX2X1 g33175(.A (wb_din_675), .B (oc5_cfg_1020), .S0 (n_8202), .Y(n_8195));
MX2X1 g33174(.A (wb_din_674), .B (n_4688), .S0 (n_8202), .Y (n_8196));
MX2X1 g33177(.A (wb_din_662), .B (n_4714), .S0 (n_8202), .Y (n_8193));
MX2X1 g33176(.A (wb_din_661), .B (oc4_cfg_1004), .S0 (n_8202), .Y(n_8194));
MX2X1 g33171(.A (wb_din_671), .B (oc5_cfg_1016), .S0 (n_8202), .Y(n_8201));
MX2X1 g33173(.A (wb_din_673), .B (n_8197), .S0 (n_8202), .Y (n_8198));
MX2X1 g33172(.A (wb_din_672), .B (n_8199), .S0 (n_8202), .Y (n_8200));
CLKBUFX1 g40977(.A (n_930), .Y (n_5732));
NAND4X1 g37086(.A (n_2445), .B (n_3398), .C (n_3404), .D (n_2244), .Y(n_5535));
MX2X1 g33179(.A (wb_din_664), .B (n_8190), .S0 (n_8202), .Y (n_8191));
MX2X1 g33178(.A (wb_din_663), .B (n_4711), .S0 (n_8202), .Y (n_8192));
INVX1 g42958(.A (u11_mem_b3_b_84 ), .Y (n_5498));
INVX2 g41112(.A (n_11852), .Y (n_4225));
AOI21X1 g37714(.A0 (n_39), .A1 (n_2553), .B0 (n_2475), .Y (n_3921));
MX2X1 g31119(.A (n_6642), .B (n_6641), .S0 (n_10267), .Y (n_10284));
MX2X1 g31118(.A (n_6496), .B (n_6495), .S0 (n_10235), .Y (n_10285));
MX2X1 g31115(.A (n_6871), .B (n_509), .S0 (n_10250), .Y (n_10289));
MX2X1 g31114(.A (n_6938), .B (n_6937), .S0 (n_10267), .Y (n_10290));
MX2X1 g31117(.A (n_6645), .B (n_6644), .S0 (n_10235), .Y (n_10287));
MX2X1 g31116(.A (n_6648), .B (n_6647), .S0 (n_10235), .Y (n_10288));
MX2X1 g31111(.A (n_6943), .B (n_6942), .S0 (n_10308), .Y (n_10295));
MX2X1 g31110(.A (n_6946), .B (n_6945), .S0 (n_10308), .Y (n_10296));
MX2X1 g31113(.A (n_6538), .B (n_6537), .S0 (n_10250), .Y (n_10291));
MX2X1 g31112(.A (n_6941), .B (n_6940), .S0 (n_10250), .Y (n_10293));
NAND2X1 g39805(.A (u7_mem_b1_b_90 ), .B (n_4225), .Y (n_4120));
INVX1 g33271(.A (n_9631), .Y (n_9672));
NAND2X1 g39803(.A (u7_mem_b2_b_59 ), .B (n_12650), .Y (n_4121));
NAND2X1 g39802(.A (n_12826), .B (u3_mem_b0_b_94 ), .Y (n_11729));
NAND2X1 g39801(.A (u7_mem_b2_b_45 ), .B (n_12641), .Y (n_4123));
NAND2X1 g39800(.A (u7_mem_b1_b_88 ), .B (n_4130), .Y (n_4124));
NAND3X1 g33276(.A (n_9579), .B (n_9472), .C (n_9471), .Y (n_9629));
NOR2X1 g40039(.A (n_2059), .B (n_2772), .Y (n_2181));
NOR2X1 g39809(.A (n_2864), .B (n_1488), .Y (n_1472));
NAND2X1 g39808(.A (u7_mem_b1_b_84 ), .B (n_4225), .Y (n_4117));
AOI22X1 g37717(.A0 (u10_din_tmp_51), .A1 (n_3339), .B0 (n_3911), .B1(in_slt_430), .Y (n_3920));
MX2X1 g38716(.A (u3_mem_b0_b_114 ), .B (wb_din_684), .S0 (n_3807), .Y(n_3627));
INVX8 g41698(.A (n_1363), .Y (n_3453));
NAND2X1 g41694(.A (n_434), .B (n_625), .Y (n_823));
INVX1 g31743(.A (n_9972), .Y (n_10344));
CLKBUFX3 g41691(.A (n_1107), .Y (n_2302));
INVX1 g41690(.A (n_2302), .Y (n_1889));
INVX1 g41693(.A (n_823), .Y (n_908));
INVX1 g41692(.A (n_823), .Y (n_1107));
INVX1 g42348(.A (u26_ps_cnt_b1_b ), .Y (n_697));
INVX1 g42349(.A (u11_mem_b3_b_65 ), .Y (n_6035));
NOR2X1 g40298(.A (n_2691), .B (n_1985), .Y (n_1979));
INVX1 g42343(.A (u10_mem_b3_b_73 ), .Y (n_6010));
INVX4 g41622(.A (n_1205), .Y (n_3543));
INVX1 g42344(.A (u10_mem_b1_b_142 ), .Y (n_1684));
INVX1 g42345(.A (u11_mem_b1_b_143 ), .Y (n_1609));
NOR2X1 g40296(.A (n_2707), .B (n_2067), .Y (n_1981));
NOR2X1 g40297(.A (n_2054), .B (n_2686), .Y (n_1980));
NAND2X1 g39135(.A (u8_mem_b2_b_32 ), .B (n_2362), .Y (n_1927));
INVX2 g41625(.A (n_909), .Y (n_1205));
NOR2X1 g40295(.A (n_2748), .B (n_1985), .Y (n_1982));
BUFX3 g41626(.A (n_909), .Y (n_1543));
NOR2X1 g40292(.A (n_2788), .B (n_2681), .Y (n_2677));
NOR2X1 g41627(.A (n_12581), .B (n_12583), .Y (n_909));
AOI21X1 g37711(.A0 (n_98), .A1 (n_2553), .B0 (n_2335), .Y (n_3922));
MX2X1 g38679(.A (u6_mem_b0_b ), .B (wb_din), .S0 (n_3632), .Y(n_3683));
NOR2X1 g40293(.A (n_2120), .B (n_2720), .Y (n_1983));
AOI21X1 g35663(.A0 (n_5906), .A1 (n_6156), .B0 (n_7120), .Y (n_7207));
NAND2X1 g39131(.A (u8_mem_b2_b_46 ), .B (n_2366), .Y (n_2352));
NOR2X1 g40291(.A (n_2780), .B (n_2686), .Y (n_2678));
AOI21X1 g35661(.A0 (n_5907), .A1 (n_5742), .B0 (n_7120), .Y (n_7117));
AOI21X1 g35660(.A0 (n_6279), .A1 (n_5760), .B0 (n_7214), .Y (n_7209));
AOI21X1 g35667(.A0 (n_5939), .A1 (n_5794), .B0 (n_7212), .Y (n_7114));
OAI21X1 g33565(.A0 (n_4413), .A1 (n_8333), .B0 (n_7992), .Y (n_8271));
AOI21X1 g35666(.A0 (n_5938), .A1 (n_5793), .B0 (n_7212), .Y (n_7172));
MX2X1 g38673(.A (u5_mem_b0_b_99 ), .B (wb_din_669), .S0 (n_3720), .Y(n_3692));
OAI21X1 g33496(.A0 (n_4863), .A1 (n_8097), .B0 (n_7575), .Y (n_8356));
AOI21X1 g35665(.A0 (n_6154), .A1 (n_6275), .B0 (n_7120), .Y (n_7204));
MX2X1 g38672(.A (u5_mem_b0_b_98 ), .B (wb_din_668), .S0 (n_841), .Y(n_3693));
AOI21X1 g35664(.A0 (n_5890), .A1 (n_6277), .B0 (n_7120), .Y (n_7205));
MX2X1 g38671(.A (u5_mem_b0_b_97 ), .B (wb_din_667), .S0 (n_3720), .Y(n_3694));
MX2X1 g38670(.A (u5_mem_b0_b_94 ), .B (wb_din_664), .S0 (n_3720), .Y(n_3696));
XOR2X1 g35722(.A (n_214), .B (n_6059), .Y (n_6060));
XOR2X1 g35723(.A (n_116), .B (n_6756), .Y (n_6757));
XOR2X1 g35721(.A (n_95), .B (n_7010), .Y (n_7011));
XOR2X1 g35726(.A (n_1446), .B (n_12588), .Y (n_6040));
MX2X1 g35727(.A (n_796), .B (u2_res_cnt_b1_b ), .S0 (n_5632), .Y(n_4843));
XOR2X1 g35724(.A (n_1255), .B (n_5964), .Y (n_5965));
XOR2X1 g35725(.A (n_1443), .B (n_5636), .Y (n_5637));
OAI21X1 g33497(.A0 (n_5121), .A1 (n_8357), .B0 (n_8075), .Y (n_8355));
MX2X1 g38675(.A (u5_mem_b0_b_95 ), .B (wb_din_665), .S0 (n_3720), .Y(n_3690));
MX2X1 g38615(.A (u4_mem_b0_b_95 ), .B (wb_din_665), .S0 (n_3765), .Y(n_3790));
MX2X1 g38674(.A (u3_mem_b0_b_95 ), .B (wb_din_665), .S0 (n_3807), .Y(n_3771));
NOR2X1 g32972(.A (n_9361), .B (n_11086), .Y (n_9516));
NOR2X1 g32973(.A (o9_empty), .B (n_12585), .Y (n_9495));
NOR2X1 g32971(.A (o8_empty), .B (n_5825), .Y (n_9496));
INVX1 g42219(.A (u10_mem_b0_b_176 ), .Y (n_1240));
NOR2X1 g32977(.A (n_9360), .B (n_11144), .Y (n_9515));
INVX1 g32974(.A (n_11126), .Y (n_9901));
AND2X1 g32975(.A (n_12502), .B (n_12636), .Y (n_11126));
NAND2X1 g32979(.A (n_8183), .B (n_8678), .Y (n_9460));
NAND2X1 g37883(.A (n_2385), .B (n_3144), .Y (n_4571));
OAI21X1 g33494(.A0 (n_4954), .A1 (n_8357), .B0 (n_8057), .Y (n_8359));
INVX1 g39114(.A (n_5282), .Y (n_4231));
INVX1 g39117(.A (n_5287), .Y (n_4230));
AOI22X1 g37330(.A0 (n_5272), .A1 (u13_intm_r_b21_b ), .B0(u13_ints_r_b21_b ), .B1 (n_4726), .Y (n_4724));
MX2X1 g38614(.A (u4_mem_b0_b_106 ), .B (wb_din_676), .S0 (n_3765), .Y(n_3791));
NAND2X1 g39110(.A (u8_mem_b2_b_54 ), .B (n_3441), .Y (n_3442));
NAND2X1 g39113(.A (u8_mem_b1_b_66 ), .B (n_12295), .Y (n_11446));
NAND2X1 g39112(.A (n_11798), .B (u8_mem_b0_b_97 ), .Y (n_11445));
AOI21X1 g38501(.A0 (u4_mem_b2_b_40 ), .A1 (n_4439), .B0 (n_2016), .Y(n_4310));
NAND2X1 g39119(.A (n_12826), .B (u3_mem_b0_b_115 ), .Y (n_3436));
NAND2X1 g39118(.A (n_3339), .B (in_slt_430), .Y (n_5287));
AOI22X1 g37336(.A0 (n_6972), .A1 (oc2_cfg_990), .B0 (u13_ints_r_b23_b), .B1 (n_3985), .Y (n_3986));
NAND2X1 g37887(.A (n_3545), .B (n_2496), .Y (n_4570));
AOI22X1 g37334(.A0 (n_5272), .A1 (u13_intm_r_b16_b ), .B0(u13_ints_r_b16_b ), .B1 (n_4726), .Y (n_4721));
OAI21X1 g33495(.A0 (n_5125), .A1 (n_8357), .B0 (n_8065), .Y (n_8358));
ADDHX1 g36200(.A (n_512), .B (n_853), .CO (n_1233), .S (n_1234));
MX2X1 g38617(.A (u7_mem_b0_b_102 ), .B (wb_din_672), .S0 (n_913), .Y(n_3786));
INVX1 g42293(.A (u26_ps_cnt_b4_b ), .Y (n_515));
ADDHX1 g36201(.A (n_606), .B (u9_wp_b2_b ), .CO (n_1557), .S (n_1558));
NAND2X1 g38859(.A (u5_mem_b3_b_140 ), .B (n_3543), .Y (n_2439));
NAND2X1 g38858(.A (u5_mem_b3_b_152 ), .B (n_3543), .Y (n_3540));
NOR2X1 g39450(.A (n_3453), .B (n_2767), .Y (n_3172));
OAI21X1 g33804(.A0 (n_3857), .A1 (n_8930), .B0 (n_8130), .Y (n_9068));
AOI21X1 g38508(.A0 (u7_mem_b3_b_131 ), .A1 (n_5145), .B0 (n_3311), .Y(n_4888));
MX2X1 g38616(.A (u4_mem_b0_b_107 ), .B (wb_din_677), .S0 (n_835), .Y(n_3788));
NOR2X1 g40319(.A (n_2705), .B (n_2741), .Y (n_2670));
MX2X1 g33157(.A (wb_din_688), .B (oc3_cfg_997), .S0 (n_8538), .Y(n_8540));
NOR2X1 g40313(.A (n_1226), .B (n_2801), .Y (n_2671));
NAND2X1 g39968(.A (u8_mem_b1_b_68 ), .B (n_12301), .Y (n_2846));
NOR2X1 g40311(.A (n_2770), .B (n_2782), .Y (n_2672));
NOR2X1 g40310(.A (n_2477), .B (n_2818), .Y (n_1969));
NOR2X1 g40317(.A (n_2059), .B (n_2732), .Y (n_1964));
NOR2X1 g40316(.A (n_2716), .B (n_2067), .Y (n_1965));
NOR2X1 g40315(.A (n_2829), .B (n_1985), .Y (n_1966));
NAND2X1 g39969(.A (u3_mem_b2_b_54 ), .B (n_3330), .Y (n_2844));
OAI21X1 g35925(.A0 (n_5682), .A1 (n_7077), .B0 (n_6191), .Y (n_7073));
MX2X1 g35996(.A (n_6647), .B (n_6646), .S0 (n_930), .Y (n_6648));
MX2X1 g38702(.A (u7_mem_b0_b_103 ), .B (wb_din_673), .S0 (n_3622), .Y(n_3647));
MX2X1 g38611(.A (u4_mem_b0_b_104 ), .B (wb_din_674), .S0 (n_3765), .Y(n_3796));
NAND2X1 g39964(.A (u4_mem_b2_b_34 ), .B (n_12079), .Y (n_2849));
NAND2X1 g39965(.A (u3_mem_b1_b_69 ), .B (n_12753), .Y (n_11720));
MX2X1 g38610(.A (u4_mem_b0_b_103 ), .B (wb_din_673), .S0 (n_3765), .Y(n_3797));
INVX1 g42321(.A (u11_mem_b1_b_133 ), .Y (n_6503));
MX2X1 g38613(.A (u7_mem_b0_b_106 ), .B (wb_din_676), .S0 (n_3622), .Y(n_3792));
OR2X1 g29969(.A (u13_ints_r_b11_b ), .B (oc3_int_set), .Y (n_10967));
OAI21X1 g33800(.A0 (n_4340), .A1 (n_8898), .B0 (n_7588), .Y (n_9072));
MX2X1 g38612(.A (u4_mem_b0_b_105 ), .B (wb_din_675), .S0 (n_3765), .Y(n_3795));
AOI22X1 g37618(.A0 (n_6641), .A1 (n_1835), .B0 (n_6450), .B1(n_1760), .Y (n_1761));
NAND2X1 g37619(.A (n_2460), .B (n_2638), .Y (n_4628));
AOI22X1 g37952(.A0 (n_2502), .A1 (n_6392), .B0 (n_6534), .B1(n_1859), .Y (n_1860));
AOI21X1 g37610(.A0 (n_6087), .A1 (n_1760), .B0 (n_1222), .Y (n_1834));
NAND2X1 g37611(.A (n_2421), .B (n_3494), .Y (n_4629));
AOI22X1 g37612(.A0 (n_2502), .A1 (n_6868), .B0 (n_6956), .B1(n_1859), .Y (n_1770));
AOI21X1 g37613(.A0 (n_6924), .A1 (n_1760), .B0 (n_1220), .Y (n_1768));
AOI22X1 g37614(.A0 (n_2502), .A1 (n_349), .B0 (n_1766), .B1 (n_1835),.Y (n_1767));
AOI22X1 g37615(.A0 (n_2502), .A1 (n_6402), .B0 (n_6551), .B1(n_1859), .Y (n_1765));
AOI22X1 g37616(.A0 (n_6644), .A1 (n_1835), .B0 (n_6617), .B1(n_1760), .Y (n_1764));
AOI22X1 g37617(.A0 (n_6495), .A1 (n_1835), .B0 (n_6614), .B1(n_1760), .Y (n_1763));
OAI21X1 g33768(.A0 (n_4928), .A1 (n_9110), .B0 (n_7760), .Y (n_9112));
OAI21X1 g33769(.A0 (n_4927), .A1 (n_9110), .B0 (n_7759), .Y (n_9111));
OAI21X1 g33760(.A0 (n_4398), .A1 (n_9110), .B0 (n_7768), .Y (n_9120));
OAI21X1 g33761(.A0 (n_4330), .A1 (n_9161), .B0 (n_7767), .Y (n_9119));
OAI21X1 g33762(.A0 (n_4457), .A1 (n_9170), .B0 (n_7766), .Y (n_9118));
OAI21X1 g33763(.A0 (n_4401), .A1 (n_9077), .B0 (n_7765), .Y (n_9117));
OAI21X1 g33764(.A0 (n_4403), .A1 (n_9077), .B0 (n_7764), .Y (n_9116));
OAI21X1 g33765(.A0 (n_4405), .A1 (n_9139), .B0 (n_7763), .Y (n_9115));
OAI21X1 g33766(.A0 (n_4415), .A1 (n_9139), .B0 (n_7762), .Y (n_9114));
OAI21X1 g33767(.A0 (n_4322), .A1 (n_9182), .B0 (n_7761), .Y (n_9113));
AOI21X1 g38413(.A0 (u8_mem_b3_b_123 ), .A1 (n_3879), .B0 (n_1495), .Y(n_3855));
NAND2X1 g37474(.A (n_4726), .B (n_5225), .Y (n_2577));
NAND2X1 g37475(.A (n_5480), .B (n_2918), .Y (n_4677));
NAND2X1 g37470(.A (u13_ints_r_b14_b ), .B (n_3985), .Y (n_2614));
BUFX3 g40860(.A (n_935), .Y (n_4439));
INVX1 g40863(.A (n_1019), .Y (n_2099));
INVX1 g40862(.A (n_1019), .Y (n_2169));
AOI21X1 g34904(.A0 (n_4845), .A1 (n_2368), .B0 (n_4805), .Y (n_6056));
NAND2X1 g37950(.A (n_2938), .B (n_3406), .Y (n_5189));
INVX4 g41193(.A (n_970), .Y (n_1406));
INVX2 g41197(.A (n_837), .Y (n_6816));
NAND2X1 g41194(.A (ic0_cfg_1026), .B (n_836), .Y (n_970));
OR2X1 g41198(.A (oc3_cfg_995), .B (n_471), .Y (n_837));
MX2X1 g34907(.A (n_4101), .B (u2_res_cnt_b3_b ), .S0 (n_5632), .Y(n_5633));
INVX1 g41874(.A (u9_mem_b3_b_62 ), .Y (n_6886));
INVX1 g42647(.A (n_445), .Y (n_765));
INVX1 g42646(.A (n_765), .Y (n_868));
INVX1 g42643(.A (u11_mem_b2_b_93 ), .Y (n_6434));
INVX1 g42642(.A (u9_mem_b0_b_170 ), .Y (n_1680));
OR2X1 g34901(.A (n_7378), .B (n_11888), .Y (n_7446));
INVX2 g42648(.A (u4_rp_b2_b ), .Y (n_445));
NAND2X1 g31612(.A (n_346), .B (n_10045), .Y (n_10035));
NAND2X1 g31613(.A (n_345), .B (n_10054), .Y (n_10034));
NAND2X1 g31610(.A (n_347), .B (n_10045), .Y (n_10038));
NAND2X1 g31611(.A (n_365), .B (n_10045), .Y (n_10037));
NAND2X1 g31616(.A (n_343), .B (n_10045), .Y (n_10030));
NAND2X1 g31617(.A (n_6089), .B (n_10045), .Y (n_10029));
NAND2X1 g31614(.A (n_2499), .B (n_10054), .Y (n_10032));
NAND2X1 g31615(.A (n_385), .B (n_10054), .Y (n_10031));
NAND2X1 g45691(.A (n_445), .B (n_551), .Y (n_12383));
INVX2 g45690(.A (n_12383), .Y (n_12384));
NAND2X1 g31618(.A (n_6087), .B (n_10073), .Y (n_10028));
NAND2X1 g31619(.A (n_5294), .B (n_10024), .Y (n_10027));
OR2X1 g34900(.A (n_7379), .B (n_11887), .Y (n_7448));
NAND2X1 g39478(.A (n_12204), .B (u6_mem_b0_b_95 ), .Y (n_11711));
INVX8 g35119(.A (n_7870), .Y (n_7496));
NOR2X1 g39477(.A (n_3117), .B (n_2786), .Y (n_3154));
OR2X1 g39475(.A (n_12640), .B (n_12634), .Y (n_1798));
NAND2X1 g39472(.A (n_12389), .B (u4_mem_b0_b_95 ), .Y (n_11666));
NAND2X1 g39473(.A (n_2344), .B (in_slt_425), .Y (n_1796));
NAND2X1 g39470(.A (u8_mem_b1_b_88 ), .B (n_12291), .Y (n_3158));
NAND2X1 g39471(.A (n_2344), .B (in_slt_431), .Y (n_1795));
OAI21X1 g36705(.A0 (n_5181), .A1 (n_5180), .B0 (n_634), .Y (n_5749));
NAND2X1 g36704(.A (n_5535), .B (n_6152), .Y (n_6093));
OAI21X1 g36707(.A0 (n_5177), .A1 (n_5176), .B0 (n_6152), .Y (n_5747));
OAI21X1 g36706(.A0 (n_4628), .A1 (n_5178), .B0 (n_6152), .Y (n_5748));
OAI21X1 g36700(.A0 (n_5179), .A1 (n_5195), .B0 (n_634), .Y (n_5753));
OAI21X1 g36702(.A0 (n_5452), .A1 (n_5453), .B0 (n_6118), .Y (n_6094));
OAI21X1 g36709(.A0 (n_4552), .A1 (n_5175), .B0 (n_6152), .Y (n_5744));
OAI21X1 g36708(.A0 (n_5174), .A1 (n_5182), .B0 (n_6152), .Y (n_5745));
INVX1 g45344(.A (n_11563), .Y (n_11564));
NAND2X1 g38851(.A (u3_mem_b3_b_142 ), .B (n_2463), .Y (n_2441));
INVX1 g39619(.A (n_5307), .Y (n_4106));
NAND2X1 g39613(.A (n_12204), .B (u6_mem_b0_b_119 ), .Y (n_3057));
NAND2X1 g39610(.A (in_slt_406), .B (n_2368), .Y (n_4776));
NAND2X1 g39611(.A (u3_mem_b1_b_63 ), .B (n_12753), .Y (n_11730));
NAND2X1 g39616(.A (n_4560), .B (in_slt_459), .Y (n_5300));
NAND2X1 g39617(.A (n_12369), .B (u6_mem_b0_b_107 ), .Y (n_3056));
NAND2X1 g39614(.A (u6_mem_b2_b_32 ), .B (n_2285), .Y (n_2276));
INVX1 g39615(.A (n_5300), .Y (n_4161));
NAND2X1 g38850(.A (u5_mem_b3_b_135 ), .B (n_1543), .Y (n_1541));
NOR2X1 g37577(.A (n_4755), .B (n_5371), .Y (n_3947));
OAI21X1 g36685(.A0 (n_4572), .A1 (n_5198), .B0 (n_784), .Y (n_6103));
NAND2X1 g38856(.A (u5_mem_b3_b_151 ), .B (n_3543), .Y (n_3542));
NOR2X1 g36415(.A (n_3432), .B (n_4837), .Y (n_4838));
OAI21X1 g33968(.A0 (n_5116), .A1 (n_8856), .B0 (n_7565), .Y (n_8857));
NAND2X1 g34649(.A (u6_mem_b2_b_52 ), .B (n_7758), .Y (n_7776));
OAI21X1 g33966(.A0 (n_4326), .A1 (n_8453), .B0 (n_7697), .Y (n_8859));
OAI21X1 g33967(.A0 (n_4321), .A1 (n_8449), .B0 (n_7566), .Y (n_8858));
OAI21X1 g33964(.A0 (n_4271), .A1 (n_8453), .B0 (n_7567), .Y (n_8861));
OAI21X1 g33965(.A0 (n_4857), .A1 (n_8097), .B0 (n_7694), .Y (n_8860));
OAI21X1 g33962(.A0 (n_4390), .A1 (n_8453), .B0 (n_7569), .Y (n_8864));
NAND2X1 g34643(.A (u6_mem_b2_b_47 ), .B (n_7758), .Y (n_7782));
NAND2X1 g34640(.A (u6_mem_b2_b_44 ), .B (n_7758), .Y (n_7785));
NAND2X1 g34641(.A (u6_mem_b2_b_45 ), .B (n_7758), .Y (n_7784));
MX2X1 g38754(.A (u8_mem_b0_b_95 ), .B (wb_din_665), .S0 (n_3826), .Y(n_3583));
NAND2X1 g38855(.A (u5_mem_b3_b_138 ), .B (n_1543), .Y (n_1336));
NOR2X1 g36414(.A (n_2577), .B (n_4837), .Y (n_4839));
MX2X1 g38755(.A (u3_mem_b0_b_119 ), .B (wb_din_689), .S0 (n_3807), .Y(n_3582));
NAND2X1 g38854(.A (u5_mem_b3_b_149 ), .B (n_3543), .Y (n_3544));
NAND2X1 g34398(.A (u4_mem_b2_b_29 ), .B (n_7984), .Y (n_8007));
NAND2X1 g34399(.A (u4_mem_b2_b_48 ), .B (n_7984), .Y (n_8006));
NAND2X1 g34468(.A (u4_mem_b3_b_127 ), .B (n_7984), .Y (n_7953));
NAND2X1 g34469(.A (u4_mem_b3_b_128 ), .B (n_7984), .Y (n_7952));
NAND2X1 g34462(.A (u4_mem_b3_b_151 ), .B (n_7984), .Y (n_7959));
NAND2X1 g34463(.A (u4_mem_b3_b_152 ), .B (n_7984), .Y (n_7958));
NAND2X1 g34460(.A (u4_mem_b3_b_150 ), .B (n_7984), .Y (n_7961));
NAND2X1 g34461(.A (u4_mem_b3_b_123 ), .B (n_7984), .Y (n_7960));
NAND2X1 g34394(.A (u4_mem_b2_b_44 ), .B (n_7984), .Y (n_8011));
NAND2X1 g34467(.A (u4_mem_b3_b_126 ), .B (n_7984), .Y (n_7954));
NAND2X1 g34464(.A (u3_mem_b1_b_70 ), .B (n_8101), .Y (n_7957));
NAND2X1 g34397(.A (u4_mem_b2_b_47 ), .B (n_7984), .Y (n_8008));
OAI21X1 g45534(.A0 (n_12146), .A1 (n_12147), .B0 (n_12149), .Y(n_12150));
MX2X1 g38756(.A (u8_mem_b0_b_99 ), .B (wb_din_669), .S0 (n_3826), .Y(n_3580));
AOI21X1 g45535(.A0 (n_12142), .A1 (n_12143), .B0 (n_12145), .Y(n_12146));
NOR2X1 g36416(.A (n_2599), .B (n_1814), .Y (n_4086));
NAND2X1 g45536(.A (n_6790), .B (u4_rp_b0_b ), .Y (n_12142));
MX2X1 g38651(.A (u5_mem_b0_b_106 ), .B (wb_din_676), .S0 (n_3720), .Y(n_3731));
NAND2X1 g45537(.A (n_145), .B (n_6803), .Y (n_12143));
NAND2X1 g36411(.A (n_6765), .B (n_6816), .Y (n_6817));
MX2X1 g38650(.A (u5_mem_b0_b_105 ), .B (wb_din_675), .S0 (n_3720), .Y(n_3732));
MX2X1 g38750(.A (u8_mem_b0_b_119 ), .B (wb_din_689), .S0 (n_3826), .Y(n_3587));
INVX1 g45538(.A (n_12144), .Y (n_12145));
MX2X1 g38653(.A (u5_mem_b0_b_108 ), .B (wb_din_678), .S0 (n_3720), .Y(n_3727));
MX2X1 g38751(.A (u3_mem_b0_b_116 ), .B (wb_din_686), .S0 (n_3807), .Y(n_3586));
MX2X1 g38652(.A (u5_mem_b0_b_107 ), .B (wb_din_677), .S0 (n_3720), .Y(n_3728));
NOR2X1 g40179(.A (n_2059), .B (n_2755), .Y (n_2060));
MX2X1 g38752(.A (u3_mem_b0_b_117 ), .B (wb_din_687), .S0 (n_3807), .Y(n_3585));
NAND2X1 g32709(.A (n_182), .B (n_10617), .Y (n_12194));
NAND3X1 g35335(.A (n_6837), .B (n_6040), .C (n_2300), .Y (n_7281));
NAND2X1 g41256(.A (n_462), .B (n_836), .Y (n_840));
NAND2X1 g36412(.A (n_6266), .B (n_12531), .Y (n_6267));
NOR2X1 g35334(.A (n_7356), .B (n_1124), .Y (n_7395));
OAI21X1 g32701(.A0 (n_5434), .A1 (n_8208), .B0 (n_8207), .Y (n_8209));
NAND2X1 g32700(.A (n_228), .B (n_10617), .Y (n_10621));
NAND2X1 g32702(.A (n_237), .B (n_10617), .Y (n_10620));
NAND2X1 g32705(.A (n_86), .B (n_10617), .Y (n_10616));
NAND2X1 g32704(.A (n_240), .B (n_10617), .Y (n_10618));
AOI21X1 g32707(.A0 (n_6205), .A1 (n_6203), .B0 (n_10617), .Y(n_10614));
NAND2X1 g32706(.A (n_328), .B (n_10617), .Y (n_10615));
AOI21X1 g38431(.A0 (u6_mem_b2_b_51 ), .A1 (n_4504), .B0 (n_2155), .Y(n_4334));
AOI21X1 g38430(.A0 (u7_mem_b1_b_72 ), .A1 (n_5118), .B0 (n_2812), .Y(n_4929));
AOI21X1 g38433(.A0 (u6_mem_b2_b_53 ), .A1 (n_4504), .B0 (n_1959), .Y(n_4332));
NOR2X1 g35440(.A (n_7025), .B (n_1271), .Y (n_7026));
AOI21X1 g38435(.A0 (u6_mem_b2_b_31 ), .A1 (n_4544), .B0 (n_1937), .Y(n_4330));
AOI21X1 g38434(.A0 (u8_mem_b2_b_39 ), .A1 (n_4499), .B0 (n_2143), .Y(n_4331));
AOI21X1 g38437(.A0 (u6_mem_b3_b ), .A1 (n_5059), .B0 (n_2964), .Y(n_4928));
AOI21X1 g38436(.A0 (u8_mem_b1_b_69 ), .A1 (n_4502), .B0 (n_2124), .Y(n_4329));
AOI21X1 g38439(.A0 (u6_mem_b3_b_132 ), .A1 (n_5059), .B0 (n_3040), .Y(n_4926));
NAND3X1 g35331(.A (n_6840), .B (n_6060), .C (n_2232), .Y (n_7282));
MX2X1 g38753(.A (u3_mem_b0_b_118 ), .B (wb_din_688), .S0 (n_3807), .Y(n_3584));
NAND3X1 g35330(.A (n_6843), .B (n_5637), .C (n_1798), .Y (n_12837));
INVX1 g35333(.A (n_7395), .Y (n_7536));
MX2X1 g38654(.A (u5_mem_b0_b_109 ), .B (wb_din_679), .S0 (n_3720), .Y(n_3725));
NAND2X1 g35444(.A (n_7303), .B (n_6673), .Y (n_7457));
INVX4 g41477(.A (n_615), .Y (n_4996));
INVX1 g41970(.A (u11_mem_b2_b_107 ), .Y (n_81));
NAND2X1 g35449(.A (n_7296), .B (n_6737), .Y (n_7452));
NAND2X1 g35448(.A (n_7299), .B (n_6693), .Y (n_7453));
MX2X1 g38657(.A (u5_mem_b0_b_111 ), .B (wb_din_681), .S0 (n_3720), .Y(n_3719));
NOR2X1 g40109(.A (n_867), .B (n_3008), .Y (n_2126));
NOR2X1 g40106(.A (n_2169), .B (n_2716), .Y (n_2129));
NOR2X1 g40107(.A (n_2761), .B (n_2864), .Y (n_2762));
NOR2X1 g40105(.A (n_2689), .B (n_2763), .Y (n_2764));
NOR2X1 g40102(.A (n_2041), .B (n_2744), .Y (n_2132));
NOR2X1 g40103(.A (n_2096), .B (n_2804), .Y (n_2131));
NOR2X1 g40100(.A (n_2133), .B (n_2794), .Y (n_2134));
NOR2X1 g40101(.A (n_2744), .B (n_2008), .Y (n_1920));
MX2X1 g37289(.A (u11_mem_b1_b_147 ), .B (n_5298), .S0 (n_6502), .Y(n_5325));
MX2X1 g37288(.A (u11_mem_b1_b_144 ), .B (n_5309), .S0 (n_6502), .Y(n_5326));
AOI21X1 g37283(.A0 (n_5333), .A1 (n_5371), .B0 (n_3948), .Y (n_5334));
MX2X1 g37282(.A (u11_mem_b1_b_138 ), .B (n_5335), .S0 (n_5405), .Y(n_5336));
MX2X1 g37281(.A (u11_mem_b2_b_107 ), .B (n_5335), .S0 (n_5312), .Y(n_5337));
MX2X1 g37280(.A (u11_mem_b1_b_148 ), .B (n_5296), .S0 (n_5405), .Y(n_5338));
MX2X1 g37287(.A (u11_mem_b1_b_142 ), .B (n_5321), .S0 (n_6502), .Y(n_5327));
MX2X1 g37286(.A (u11_mem_b1_b_141 ), .B (n_5313), .S0 (n_6502), .Y(n_5329));
MX2X1 g37285(.A (u10_mem_b2_b_117 ), .B (n_5330), .S0 (n_5341), .Y(n_5331));
MX2X1 g37284(.A (u11_mem_b1_b_140 ), .B (n_5315), .S0 (n_6502), .Y(n_5332));
MX2X1 g38656(.A (u5_mem_b0_b_110 ), .B (wb_din_680), .S0 (n_3720), .Y(n_3722));
AOI21X1 g38158(.A0 (u4_mem_b2_b_49 ), .A1 (n_4439), .B0 (n_1992), .Y(n_4428));
AOI21X1 g38404(.A0 (u6_mem_b1_b ), .A1 (n_5112), .B0 (n_2675), .Y(n_4948));
INVX1 g42784(.A (ic2_cfg_1049), .Y (n_518));
AOI21X1 g38405(.A0 (u6_mem_b1_b_70 ), .A1 (n_5112), .B0 (n_2652), .Y(n_4947));
INVX1 g42785(.A (u11_mem_b1_b_137 ), .Y (n_1644));
AOI21X1 g38406(.A0 (u7_mem_b2_b_32 ), .A1 (n_4540), .B0 (n_2204), .Y(n_4339));
MX2X1 g38738(.A (u8_mem_b0_b_100 ), .B (wb_din_670), .S0 (n_3826), .Y(n_3602));
MX2X1 g38659(.A (u5_mem_b0_b_113 ), .B (wb_din_683), .S0 (n_3720), .Y(n_3715));
AOI21X1 g38155(.A0 (u4_mem_b2_b_47 ), .A1 (n_4439), .B0 (n_1969), .Y(n_4430));
AOI21X1 g38400(.A0 (u8_mem_b1_b_65 ), .A1 (n_4502), .B0 (n_2193), .Y(n_4340));
INVX1 g36979(.A (n_6779), .Y (n_6075));
AOI21X1 g38401(.A0 (u5_mem_b3_b_127 ), .A1 (n_4996), .B0 (n_3031), .Y(n_4950));
NAND4X1 g36976(.A (n_11715), .B (n_11716), .C (n_1810), .D (n_2426),.Y (n_5833));
XOR2X1 g38402(.A (u9_rp_b2_b ), .B (n_737), .Y (n_1085));
OAI21X1 g35949(.A0 (n_5529), .A1 (n_7063), .B0 (n_5896), .Y (n_6977));
AOI21X1 g38403(.A0 (u7_mem_b3_b_136 ), .A1 (n_4961), .B0 (n_3501), .Y(n_4949));
MX2X1 g38739(.A (u3_mem_b0_b_108 ), .B (wb_din_678), .S0 (n_3807), .Y(n_3601));
INVX1 g41802(.A (u9_mem_b3_b_73 ), .Y (n_6951));
MX2X1 g36065(.A (n_6881), .B (n_6920), .S0 (n_6898), .Y (n_6882));
AOI22X1 g37672(.A0 (in_slt_403), .A1 (n_1406), .B0 (u9_din_tmp_48),.B1 (n_4616), .Y (n_4614));
AOI22X1 g37673(.A0 (in_slt_406), .A1 (n_3415), .B0 (in_slt_404), .B1(n_3935), .Y (n_3932));
AOI21X1 g38374(.A0 (u8_mem_b2_b_41 ), .A1 (n_4499), .B0 (n_2292), .Y(n_4350));
AOI22X1 g37671(.A0 (n_347), .A1 (n_1835), .B0 (n_5333), .B1 (n_1760),.Y (n_1699));
AOI22X1 g37676(.A0 (n_2502), .A1 (n_6404), .B0 (n_6647), .B1(n_1835), .Y (n_1697));
MX2X1 g38736(.A (u8_mem_b0_b ), .B (wb_din), .S0 (n_3826), .Y(n_3604));
INVX1 g36995(.A (n_12368), .Y (n_5704));
AOI21X1 g38373(.A0 (u8_mem_b3_b_128 ), .A1 (n_3879), .B0 (n_1480), .Y(n_3861));
AOI22X1 g37674(.A0 (n_3415), .A1 (in_slt_407), .B0 (n_1406), .B1(in_slt_405), .Y (n_4613));
AOI22X1 g37869(.A0 (n_1756), .A1 (n_5947), .B0 (n_5984), .B1(n_1643), .Y (n_1567));
NAND2X1 g37868(.A (n_2458), .B (n_3468), .Y (n_12059));
AOI22X1 g37866(.A0 (n_6431), .A1 (n_1575), .B0 (n_6650), .B1(n_1831), .Y (n_1832));
NAND2X1 g37865(.A (n_4229), .B (n_3070), .Y (n_5203));
AOI22X1 g37675(.A0 (n_6638), .A1 (n_1835), .B0 (n_6505), .B1(n_1760), .Y (n_1698));
NAND2X1 g37863(.A (n_2388), .B (n_3480), .Y (n_4576));
AOI22X1 g37862(.A0 (n_1756), .A1 (n_6344), .B0 (n_6484), .B1(n_1643), .Y (n_1569));
AOI22X1 g37861(.A0 (u10_din_tmp_52), .A1 (n_3339), .B0 (n_3911), .B1(in_slt_431), .Y (n_3913));
NAND2X1 g37860(.A (n_4163), .B (n_3073), .Y (n_12052));
MX2X1 g33159(.A (wb_din_662), .B (oc0_cfg_965), .S0 (n_8538), .Y(n_8535));
MX2X1 g33158(.A (wb_din_689), .B (n_8536), .S0 (n_8538), .Y (n_8537));
MX2X1 g33156(.A (wb_din_687), .B (oc3_cfg_996), .S0 (n_8538), .Y(n_8542));
MX2X1 g33155(.A (wb_din_686), .B (oc3_cfg_995), .S0 (n_8538), .Y(n_8543));
MX2X1 g33154(.A (wb_din_685), .B (oc3_cfg_994), .S0 (n_8538), .Y(n_8545));
MX2X1 g33153(.A (wb_din_684), .B (n_1873), .S0 (n_8538), .Y (n_8546));
MX2X1 g33152(.A (wb_din_683), .B (oc2_cfg_990), .S0 (n_8538), .Y(n_8548));
MX2X1 g33151(.A (wb_din_682), .B (n_3987), .S0 (n_8538), .Y (n_8549));
MX2X1 g33150(.A (wb_din_681), .B (n_8550), .S0 (n_8538), .Y (n_8551));
MX2X1 g31137(.A (n_6621), .B (n_6620), .S0 (n_10747), .Y (n_10262));
MX2X1 g31136(.A (n_6926), .B (n_6924), .S0 (n_10277), .Y (n_10263));
MX2X1 g31135(.A (n_6894), .B (n_6893), .S0 (n_10277), .Y (n_10264));
MX2X1 g31134(.A (n_6629), .B (n_6628), .S0 (n_10267), .Y (n_10265));
MX2X1 g31133(.A (n_6929), .B (n_6928), .S0 (n_10267), .Y (n_10266));
MX2X1 g31132(.A (n_6624), .B (n_6623), .S0 (n_9724), .Y (n_10651));
MX2X1 g31131(.A (n_6901), .B (n_6900), .S0 (n_10267), .Y (n_10268));
MX2X1 g31139(.A (n_6615), .B (n_6614), .S0 (n_10235), .Y (n_10259));
MX2X1 g31138(.A (n_6619), .B (n_6617), .S0 (n_10747), .Y (n_10261));
MX2X1 g38734(.A (u7_mem_b0_b_117 ), .B (wb_din_687), .S0 (n_3622), .Y(n_3607));
INVX1 g42078(.A (u9_mem_b3_b_72 ), .Y (n_6922));
NOR2X1 g39861(.A (n_5059), .B (n_2691), .Y (n_2916));
NAND2X1 g39860(.A (u7_mem_b1_b_73 ), .B (n_11856), .Y (n_4113));
NAND2X1 g39863(.A (n_12721), .B (u3_mem_b0_b_103 ), .Y (n_2914));
NAND2X1 g39862(.A (u8_mem_b1_b_86 ), .B (n_12291), .Y (n_2915));
NOR2X1 g39865(.A (n_3089), .B (n_2829), .Y (n_2912));
NAND2X1 g39864(.A (u3_mem_b2_b_49 ), .B (n_3330), .Y (n_2913));
NOR2X1 g39867(.A (u11_mem_b2_b_100 ), .B (n_1214), .Y (n_1211));
NOR2X1 g39866(.A (n_2794), .B (n_1488), .Y (n_1414));
NAND2X1 g39869(.A (n_12204), .B (u6_mem_b0_b_98 ), .Y (n_11717));
INVX1 g41780(.A (n_12332), .Y (n_438));
MX2X1 g38735(.A (u3_mem_b0_b_103 ), .B (wb_din_673), .S0 (n_3807), .Y(n_3606));
OAI21X1 g33874(.A0 (n_4907), .A1 (n_8981), .B0 (n_7650), .Y (n_8980));
NAND2X1 g38991(.A (u6_mem_b3_b_124 ), .B (n_12622), .Y (n_2376));
INVX1 g41803(.A (u9_mem_b2_b_105 ), .Y (n_1766));
OAI21X1 g33870(.A0 (n_4294), .A1 (n_9010), .B0 (n_7655), .Y (n_8985));
INVX4 g33359(.A (n_9703), .Y (n_9873));
MX2X1 g38733(.A (u6_mem_b0_b_111 ), .B (wb_din_681), .S0 (n_3632), .Y(n_3608));
OR2X1 g41485_dup(.A (n_485), .B (n_422), .Y (n_12802));
NAND2X1 g38997(.A (u5_mem_b3_b_141 ), .B (n_3543), .Y (n_3526));
INVX1 g35256(.A (o8_status_1002), .Y (n_7035));
AOI22X1 g35705(.A0 (n_6686), .A1 (i6_dout_637), .B0 (i3_dout_575),.B1 (n_6700), .Y (n_6677));
INVX1 g35254(.A (o7_status_992), .Y (n_7036));
AOI22X1 g35707(.A0 (n_6686), .A1 (i6_dout_638), .B0 (i3_dout_576),.B1 (n_6700), .Y (n_6676));
INVX1 g35252(.A (o6_status_982), .Y (n_7160));
AOI22X1 g35701(.A0 (n_6686), .A1 (i6_dout_633), .B0 (i3_dout_571),.B1 (n_6700), .Y (n_6683));
INVX1 g35250(.A (o4_status_972), .Y (n_7161));
AOI22X1 g35703(.A0 (n_6686), .A1 (i6_dout_626), .B0 (i3_dout_564),.B1 (n_6700), .Y (n_6680));
NOR2X1 g40119(.A (n_2470), .B (n_2790), .Y (n_2115));
AOI22X1 g35708(.A0 (n_6686), .A1 (i6_dout_635), .B0 (i3_dout_573),.B1 (n_6700), .Y (n_6675));
AOI22X1 g35709(.A0 (n_5892), .A1 (n_7443), .B0 (u13_ints_r_b1_b ), .B1(n_3985), .Y (n_7113));
INVX1 g35258(.A (o9_status_1012), .Y (n_7034));
MX2X1 g38731(.A (u7_mem_b0_b_119 ), .B (wb_din_689), .S0 (n_3622), .Y(n_3610));
INVX1 g42365(.A (ic2_int_set_724), .Y (n_749));
INVX1 g42360(.A (in_slt_739), .Y (n_221));
INVX1 g42362(.A (n_4703), .Y (n_699));
NOR2X1 g41067(.A (n_5588), .B (n_802), .Y (n_9444));
INVX1 g43015(.A (ic1_cfg_1039), .Y (n_523));
INVX1 g43014(.A (n_523), .Y (n_4687));
INVX8 g32958(.A (n_9903), .Y (n_10820));
NOR2X1 g40110(.A (n_2691), .B (n_2067), .Y (n_2124));
NOR2X1 g39289(.A (n_3486), .B (n_2801), .Y (n_3313));
AOI22X1 g37836(.A0 (n_125), .A1 (n_1575), .B0 (n_5524), .B1 (n_1831),.Y (n_1590));
NAND2X1 g39139(.A (n_12389), .B (u4_mem_b0_b_114 ), .Y (n_2700));
NAND2X1 g39138(.A (u4_mem_b1_b_73 ), .B (n_12261), .Y (n_11472));
NOR2X1 g39136(.A (n_5138), .B (n_2765), .Y (n_3426));
NOR2X1 g40294(.A (n_2736), .B (n_2691), .Y (n_2676));
NAND2X1 g39134(.A (u4_mem_b2_b_37 ), .B (n_12079), .Y (n_2644));
NOR2X1 g39133(.A (n_3089), .B (n_2732), .Y (n_3428));
NAND2X1 g39132(.A (n_1377), .B (u6_rp_b3_b ), .Y (n_4834));
AOI22X1 g37837(.A0 (n_1756), .A1 (n_6357), .B0 (n_6498), .B1(n_1643), .Y (n_1588));
NAND2X1 g45906(.A (n_12637), .B (n_12638), .Y (n_12639));
NAND2X1 g39332(.A (u5_mem_b2_b ), .B (n_12823), .Y (n_11494));
AOI22X1 g37830(.A0 (n_1756), .A1 (n_1600), .B0 (n_1599), .B1(n_1643), .Y (n_1601));
MX2X1 g34075(.A (u6_mem_b0_b_95 ), .B (n_3664), .S0 (n_7505), .Y(n_8756));
MX2X1 g34074(.A (u6_mem_b0_b_94 ), .B (n_3648), .S0 (n_7505), .Y(n_9405));
MX2X1 g34077(.A (u6_mem_b0_b_97 ), .B (n_3663), .S0 (n_7505), .Y(n_9404));
MX2X1 g34076(.A (u6_mem_b0_b_96 ), .B (n_3652), .S0 (n_7505), .Y(n_8755));
MX2X1 g34071(.A (u6_mem_b0_b_120 ), .B (n_3667), .S0 (n_7505), .Y(n_8759));
MX2X1 g34073(.A (u6_mem_b0_b_93 ), .B (n_3628), .S0 (n_7505), .Y(n_8758));
MX2X1 g34072(.A (u6_mem_b0_b_121 ), .B (n_3666), .S0 (n_7505), .Y(n_9406));
MX2X1 g34079(.A (u6_mem_b0_b_99 ), .B (n_3658), .S0 (n_7505), .Y(n_9402));
MX2X1 g34078(.A (u6_mem_b0_b_98 ), .B (n_3660), .S0 (n_7505), .Y(n_8754));
AOI22X1 g37831(.A0 (n_1756), .A1 (n_1596), .B0 (n_1595), .B1(n_1643), .Y (n_1597));
NOR2X1 g39276(.A (u10_mem_b1_b_139 ), .B (n_2364), .Y (n_2475));
AOI22X1 g37832(.A0 (n_188), .A1 (n_1575), .B0 (n_5498), .B1 (n_1831),.Y (n_1594));
AOI22X1 g37774(.A0 (n_1756), .A1 (n_6363), .B0 (n_6466), .B1(n_1575), .Y (n_1662));
NAND2X1 g38934(.A (u7_mem_b3_b_149 ), .B (n_1546), .Y (n_1523));
AND2X1 g41730(.A (n_568), .B (n_936), .Y (n_7528));
AOI22X1 g37833(.A0 (n_1756), .A1 (n_1592), .B0 (n_1591), .B1(n_1643), .Y (n_1593));
NAND2X1 g37499(.A (n_6972), .B (n_8536), .Y (n_4665));
NOR2X1 g37497(.A (n_5292), .B (n_6594), .Y (n_4666));
NAND2X1 g38935(.A (u8_mem_b3_b_150 ), .B (n_2468), .Y (n_2400));
AOI21X1 g38376(.A0 (u7_mem_b1_b_81 ), .A1 (n_5069), .B0 (n_2793), .Y(n_4964));
AOI21X1 g38377(.A0 (u3_mem_b1_b_77 ), .A1 (n_5157), .B0 (n_2653), .Y(n_4963));
AOI22X1 g37670(.A0 (in_slt_402), .A1 (n_1406), .B0 (u9_din_tmp_47),.B1 (n_4616), .Y (n_4615));
XOR2X1 g38375(.A (n_116), .B (n_4996), .Y (n_4349));
AOI21X1 g38372(.A0 (u5_mem_b3_b_130 ), .A1 (n_4996), .B0 (n_3058), .Y(n_4965));
NAND2X1 g37677(.A (n_2374), .B (n_2863), .Y (n_4611));
AOI21X1 g38370(.A0 (u6_mem_b1_b_77 ), .A1 (n_5019), .B0 (n_2809), .Y(n_4967));
AOI21X1 g38371(.A0 (u5_mem_b3_b_129 ), .A1 (n_4996), .B0 (n_2854), .Y(n_4966));
NAND2X1 g37678(.A (n_4109), .B (n_3134), .Y (n_5224));
AOI22X1 g37679(.A0 (n_6940), .A1 (n_1859), .B0 (n_6909), .B1(n_1760), .Y (n_1696));
AOI21X1 g38378(.A0 (u8_mem_b3_b_151 ), .A1 (n_3879), .B0 (n_1472), .Y(n_3860));
AOI21X1 g38379(.A0 (u7_mem_b3_b_137 ), .A1 (n_4961), .B0 (n_3455), .Y(n_4962));
OAI21X1 g33702(.A0 (n_4346), .A1 (n_8856), .B0 (n_7835), .Y (n_9195));
OAI21X1 g33703(.A0 (n_3850), .A1 (n_8453), .B0 (n_7727), .Y (n_9193));
OAI21X1 g33700(.A0 (n_3858), .A1 (n_8464), .B0 (n_7837), .Y (n_9197));
OAI21X1 g33701(.A0 (n_4319), .A1 (n_8433), .B0 (n_7596), .Y (n_9196));
OAI21X1 g33706(.A0 (n_4947), .A1 (n_9182), .B0 (n_7830), .Y (n_9190));
OAI21X1 g33707(.A0 (n_4933), .A1 (n_9182), .B0 (n_7828), .Y (n_9189));
OAI21X1 g33704(.A0 (n_4948), .A1 (n_9161), .B0 (n_7832), .Y (n_9192));
OAI21X1 g33705(.A0 (n_4930), .A1 (n_9161), .B0 (n_7831), .Y (n_9191));
OAI21X1 g33708(.A0 (n_4946), .A1 (n_9182), .B0 (n_7827), .Y (n_9188));
OAI21X1 g33709(.A0 (n_4938), .A1 (n_9161), .B0 (n_7825), .Y (n_9187));
OAI21X1 g33957(.A0 (n_4872), .A1 (n_8911), .B0 (n_7572), .Y (n_8870));
NAND2X1 g38937(.A (u7_mem_b3_b_139 ), .B (n_1538), .Y (n_1521));
INVX1 g41898(.A (u10_mem_b3_b_79 ), .Y (n_5516));
NOR2X1 g37498(.A (n_4745), .B (n_6594), .Y (n_3959));
NOR2X1 g37496(.A (n_4769), .B (n_5371), .Y (n_3960));
OAI21X1 g33956(.A0 (n_4278), .A1 (n_8868), .B0 (n_7573), .Y (n_8871));
NOR2X1 g37495(.A (n_4772), .B (n_5371), .Y (n_3961));
NOR2X1 g37492(.A (n_4747), .B (n_5371), .Y (n_4085));
NAND2X1 g37493(.A (n_5480), .B (n_3137), .Y (n_4667));
NAND2X1 g37490(.A (n_5480), .B (n_3138), .Y (n_4669));
NAND2X1 g37491(.A (n_5480), .B (n_3275), .Y (n_4668));
NAND2X1 g38930(.A (u7_mem_b3_b_130 ), .B (n_1538), .Y (n_1526));
OAI21X1 g33955(.A0 (n_4270), .A1 (n_8891), .B0 (n_7580), .Y (n_8872));
NAND2X1 g38931(.A (u7_mem_b3_b_145 ), .B (n_1546), .Y (n_1525));
INVX8 g41278(.A (n_1055), .Y (n_3720));
OR2X1 g38932(.A (n_1484), .B (n_680), .Y (n_1104));
INVX1 g42973(.A (u10_mem_b1_b_124 ), .Y (n_6408));
INVX1 g42621(.A (u11_mem_b0_b_172 ), .Y (n_1620));
AOI22X1 g37819(.A0 (n_2558), .A1 (n_5945), .B0 (n_6021), .B1(n_2534), .Y (n_2526));
INVX1 g42990(.A (n_5825), .Y (n_1481));
INVX2 g42625(.A (u3_wp_b0_b ), .Y (n_627));
INVX4 g42624(.A (n_627), .Y (n_1424));
INVX1 g42995(.A (oc4_cfg), .Y (n_418));
CLKBUFX1 g42994(.A (n_418), .Y (n_5825));
INVX1 g42629(.A (u11_mem_b2_b_98 ), .Y (n_433));
INVX1 g42998(.A (u10_mem_b1_b_132 ), .Y (n_508));
INVX1 g40842(.A (n_1167), .Y (n_2006));
NAND4X1 g45900(.A (n_4175), .B (n_4191), .C (n_2993), .D (n_1339), .Y(n_12627));
NAND2X1 g39334(.A (u5_mem_b1_b_65 ), .B (n_3257), .Y (n_12807));
NAND2X1 g31638(.A (n_5514), .B (n_10010), .Y (n_10006));
NAND2X1 g31639(.A (n_5512), .B (n_10010), .Y (n_10005));
NAND2X2 g40844(.A (n_710), .B (u5_wp_b1_b ), .Y (n_867));
NAND2X1 g31634(.A (n_5520), .B (n_10010), .Y (n_10011));
NAND2X1 g31635(.A (n_5363), .B (n_10081), .Y (n_10009));
NAND2X1 g31636(.A (n_5518), .B (n_10010), .Y (n_10008));
NAND2X1 g31637(.A (n_5516), .B (n_10065), .Y (n_10007));
NAND3X1 g31630(.A (n_11564), .B (n_1203), .C (n_9514), .Y (n_9759));
NAND2X1 g31631(.A (n_6680), .B (n_9454), .Y (n_9608));
NAND2X1 g31632(.A (n_5577), .B (n_10081), .Y (n_10013));
NAND2X1 g31633(.A (n_5575), .B (n_10081), .Y (n_10012));
NOR2X1 g41710(.A (u13_ints_r_b15_b ), .B (n_668), .Y (n_669));
NAND2X1 g39459(.A (n_12826), .B (u3_mem_b0_b_95 ), .Y (n_11737));
INVX1 g35138(.A (n_7402), .Y (n_8981));
OAI21X1 g30949(.A0 (n_4793), .A1 (n_10450), .B0 (n_10079), .Y(n_10769));
OAI21X1 g30948(.A0 (n_5380), .A1 (n_10450), .B0 (n_10080), .Y(n_10770));
INVX8 g41717(.A (n_1106), .Y (n_3632));
OAI21X1 g30945(.A0 (n_977), .A1 (o9_status), .B0 (n_9550), .Y(n_9581));
OAI21X1 g30944(.A0 (n_847), .A1 (o8_status), .B0 (n_9552), .Y(n_9582));
OAI21X1 g30947(.A0 (n_5425), .A1 (n_10450), .B0 (n_10082), .Y(n_10771));
OAI21X1 g30946(.A0 (n_5426), .A1 (n_10679), .B0 (n_10084), .Y(n_10772));
OAI21X1 g30941(.A0 (n_1381), .A1 (o4_status), .B0 (n_9606), .Y(n_9644));
CLKBUFX1 g35136(.A (o6_we), .Y (n_7408));
INVX2 g35135(.A (n_7408), .Y (n_9286));
OAI21X1 g30942(.A0 (n_1391), .A1 (o6_status), .B0 (n_9554), .Y(n_9583));
OAI21X1 g36729(.A0 (n_2302), .A1 (n_5420), .B0 (n_4036), .Y (n_5421));
AOI21X1 g36728(.A0 (n_5575), .A1 (n_6594), .B0 (n_4819), .Y (n_5576));
AOI21X1 g36727(.A0 (n_5577), .A1 (n_6594), .B0 (n_4820), .Y (n_5578));
OAI21X1 g36726(.A0 (n_2368), .A1 (n_4074), .B0 (n_1813), .Y (n_4075));
AOI21X1 g36725(.A0 (n_6087), .A1 (n_5371), .B0 (n_5569), .Y (n_6088));
AOI21X1 g36724(.A0 (n_6089), .A1 (n_5371), .B0 (n_5570), .Y (n_6090));
MX2X1 g36723(.A (u9_mem_b2_b_106 ), .B (n_5733), .S0 (n_5732), .Y(n_5734));
MX2X1 g36722(.A (u9_mem_b2_b_105 ), .B (n_5736), .S0 (n_5732), .Y(n_5735));
MX2X1 g36721(.A (u10_mem_b1_b_137 ), .B (n_5422), .S0 (n_5407), .Y(n_5423));
MX2X1 g36720(.A (u9_mem_b1_b_136 ), .B (n_5736), .S0 (n_5730), .Y(n_5737));
INVX1 g42199(.A (n_625), .Y (n_4690));
OR2X1 g32978_dup(.A (n_9717), .B (n_9666), .Y (n_11894));
INVX1 g42191(.A (n_760), .Y (n_680));
INVX1 g42197(.A (u9_mem_b2_b_114 ), .Y (n_346));
INVX1 g42166(.A (u9_mem_b1_b_133 ), .Y (n_6528));
INVX1 g42195(.A (u11_mem_b2_b_113 ), .Y (n_298));
INVX1 g42194(.A (u11_mem_b3_b_63 ), .Y (n_6625));
OAI21X1 g33950(.A0 (n_4495), .A1 (n_8438), .B0 (n_7577), .Y (n_8879));
NAND2X1 g34310(.A (u3_mem_b3_b_146 ), .B (n_8101), .Y (n_8086));
INVX1 g41520(.A (n_1122), .Y (n_1379));
OAI21X1 g33471(.A0 (n_4873), .A1 (n_8387), .B0 (n_8102), .Y (n_8388));
NAND2X1 g34312(.A (u3_mem_b3_b_148 ), .B (n_8141), .Y (n_8084));
MX2X1 g38770(.A (u6_mem_b0_b_101 ), .B (wb_din_671), .S0 (n_813), .Y(n_3565));
NAND2X1 g34313(.A (u3_mem_b3_b_149 ), .B (n_8101), .Y (n_8083));
NAND2X1 g34314(.A (u3_mem_b3_b_150 ), .B (n_8101), .Y (n_8081));
NAND2X1 g34315(.A (u3_mem_b3_b_123 ), .B (n_8141), .Y (n_8082));
MX2X1 g31090(.A (n_6665), .B (n_6664), .S0 (n_10137), .Y (n_10321));
MX2X1 g31091(.A (n_6663), .B (n_6662), .S0 (n_10315), .Y (n_10319));
MX2X1 g31092(.A (n_6661), .B (n_6660), .S0 (n_10137), .Y (n_10318));
MX2X1 g31093(.A (n_6034), .B (n_6033), .S0 (n_10315), .Y (n_10317));
MX2X1 g31094(.A (n_6031), .B (n_6030), .S0 (n_10315), .Y (n_10316));
OAI21X1 g33476(.A0 (n_5137), .A1 (n_8380), .B0 (n_8095), .Y (n_8381));
MX2X1 g31096(.A (n_6957), .B (n_6956), .S0 (n_10235), .Y (n_10314));
MX2X1 g31097(.A (n_6657), .B (n_6656), .S0 (n_10235), .Y (n_10313));
MX2X1 g31098(.A (n_6552), .B (n_6551), .S0 (n_10267), .Y (n_10311));
MX2X1 g31099(.A (n_6541), .B (n_6540), .S0 (n_10308), .Y (n_10310));
NAND2X1 g34317(.A (u8_mem_b3_b_149 ), .B (n_7976), .Y (n_8080));
NAND2X1 g34318(.A (u3_mem_b3_b_152 ), .B (n_8141), .Y (n_8079));
NAND2X1 g34319(.A (u7_mem_b2_b_29 ), .B (n_7651), .Y (n_8078));
NAND2X1 g38938(.A (u7_mem_b3_b_122 ), .B (n_1538), .Y (n_1362));
INVX1 g42626(.A (u10_mem_b3_b_86 ), .Y (n_5506));
NAND2X1 g34668(.A (u6_mem_b3_b_133 ), .B (n_7758), .Y (n_7756));
OAI21X1 g33949(.A0 (n_4864), .A1 (n_8911), .B0 (n_7578), .Y (n_8880));
OAI21X1 g33940(.A0 (n_4866), .A1 (n_8856), .B0 (n_7585), .Y (n_8893));
OAI21X1 g33941(.A0 (n_4328), .A1 (n_8891), .B0 (n_7584), .Y (n_8892));
OAI21X1 g33942(.A0 (n_4273), .A1 (n_8433), .B0 (n_7583), .Y (n_8890));
OAI21X1 g33943(.A0 (n_4865), .A1 (n_8856), .B0 (n_7791), .Y (n_8888));
NAND2X1 g34664(.A (u6_mem_b2_b_37 ), .B (n_7758), .Y (n_7761));
NAND2X1 g34665(.A (u6_mem_b3_b ), .B (n_7758), .Y (n_7760));
OAI21X1 g33946(.A0 (n_4963), .A1 (n_8440), .B0 (n_7581), .Y (n_8883));
OAI21X1 g33947(.A0 (n_4350), .A1 (n_8433), .B0 (n_8125), .Y (n_8882));
NAND2X1 g38939(.A (u4_mem_b3_b_144 ), .B (n_3556), .Y (n_3530));
NAND2X1 g34761(.A (u7_mem_b2_b_48 ), .B (n_7651), .Y (n_7673));
NAND2X1 g39634(.A (n_2325), .B (in_slt6), .Y (n_2273));
NAND2X1 g39635(.A (u4_mem_b1_b_87 ), .B (n_12267), .Y (n_4155));
NAND2X1 g39636(.A (u6_mem_b2_b_33 ), .B (n_2285), .Y (n_2272));
NAND2X1 g39637(.A (u3_mem_b1_b_88 ), .B (n_3316), .Y (n_3045));
NAND2X1 g39630(.A (u6_mem_b2_b_29 ), .B (n_3474), .Y (n_12819));
NAND2X1 g39631(.A (u5_mem_b1_b_60 ), .B (n_3236), .Y (n_11442));
NAND2X1 g39632(.A (u6_mem_b1_b_62 ), .B (n_12169), .Y (n_12822));
NAND2X1 g39633(.A (u6_mem_b2_b_31 ), .B (n_3474), .Y (n_12821));
NAND2X1 g39638(.A (n_3252), .B (u7_mem_b0_b_114 ), .Y (n_3044));
NAND2X1 g39639(.A (n_3259), .B (u5_mem_b0_b_121 ), .Y (n_3043));
OAI21X1 g33492(.A0 (n_5130), .A1 (n_8375), .B0 (n_7619), .Y (n_8361));
OAI21X1 g33493(.A0 (n_4953), .A1 (n_8375), .B0 (n_8079), .Y (n_8360));
NAND2X1 g34440(.A (u4_mem_b3_b_138 ), .B (n_7984), .Y (n_7974));
NAND2X1 g34441(.A (u4_mem_b3_b_139 ), .B (n_7984), .Y (n_7973));
NAND2X1 g34442(.A (u4_mem_b3_b_140 ), .B (n_7984), .Y (n_7972));
NAND2X1 g34443(.A (u4_mem_b3_b_122 ), .B (n_7984), .Y (n_7971));
NOR2X1 g41413(.A (n_680), .B (n_515), .Y (n_681));
OAI21X1 g33498(.A0 (n_5124), .A1 (n_8357), .B0 (n_8074), .Y (n_8354));
OAI21X1 g33499(.A0 (n_4908), .A1 (n_8387), .B0 (n_8073), .Y (n_8353));
INVX2 g34449(.A (n_7515), .Y (n_8611));
INVX1 g34919(.A (n_7428), .Y (n_9110));
AOI21X1 g45516(.A0 (n_12120), .A1 (n_12121), .B0 (n_12640), .Y(n_12124));
AOI21X1 g38446(.A0 (u6_mem_b3_b_142 ), .A1 (n_5100), .B0 (n_3167), .Y(n_4921));
INVX1 g42256(.A (u10_mem_b2_b_92 ), .Y (n_6623));
INVX1 g42525(.A (u11_mem_b1_b_135 ), .Y (n_5988));
ADDHX1 g38778(.A (u2_to_cnt_b0_b ), .B (u2_to_cnt_b1_b ), .CO (n_1553),.S (n_795));
INVX1 g42253(.A (u9_mem_b2_b_106 ), .Y (n_141));
NAND2X1 g32723(.A (n_109), .B (n_10605), .Y (n_11748));
NAND2X1 g32722(.A (n_281), .B (n_10605), .Y (n_12453));
NAND2X1 g32721(.A (n_282), .B (n_10605), .Y (n_10599));
NAND2X1 g32720(.A (n_267), .B (n_10605), .Y (n_10601));
NAND2X1 g32727(.A (n_329), .B (n_10605), .Y (n_10592));
NAND2X1 g32726(.A (n_308), .B (n_10583), .Y (n_11634));
NAND2X1 g32725(.A (n_9873), .B (n_8182), .Y (n_11096));
NAND2X1 g32724(.A (n_16), .B (n_10605), .Y (n_10595));
NAND2X1 g32729(.A (n_152), .B (n_10583), .Y (n_11616));
NAND2X1 g32728(.A (n_302), .B (n_10583), .Y (n_11614));
OR2X1 g45453(.A (n_9719), .B (n_9668), .Y (n_11891));
OR2X1 g45452(.A (n_12636), .B (n_12501), .Y (n_11889));
MX2X1 g38636(.A (u4_mem_b0_b_96 ), .B (wb_din_666), .S0 (n_3765), .Y(n_3755));
INVX1 g45451(.A (n_11852), .Y (n_11856));
AOI21X1 g38419(.A0 (u6_mem_b1_b_62 ), .A1 (n_5019), .B0 (n_2811), .Y(n_4935));
AOI21X1 g38418(.A0 (u6_mem_b1_b_90 ), .A1 (n_5019), .B0 (n_2750), .Y(n_4936));
AOI21X1 g38149(.A0 (u8_mem_b2_b_56 ), .A1 (n_4491), .B0 (n_1989), .Y(n_4434));
AOI21X1 g38148(.A0 (u4_mem_b2_b_43 ), .A1 (n_4439), .B0 (n_2188), .Y(n_4435));
AOI21X1 g38145(.A0 (u4_mem_b2_b_39 ), .A1 (n_4439), .B0 (n_2129), .Y(n_4440));
AOI21X1 g38411(.A0 (u6_mem_b1_b_79 ), .A1 (n_5019), .B0 (n_2664), .Y(n_4942));
AOI21X1 g38410(.A0 (u6_mem_b1_b_60 ), .A1 (n_5019), .B0 (n_2709), .Y(n_4943));
AOI21X1 g38417(.A0 (u6_mem_b1_b_61 ), .A1 (n_5019), .B0 (n_2824), .Y(n_4937));
AOI21X1 g38416(.A0 (u6_mem_b1_b_73 ), .A1 (n_5019), .B0 (n_2680), .Y(n_4938));
AOI21X1 g38415(.A0 (u6_mem_b1_b_87 ), .A1 (n_5019), .B0 (n_2826), .Y(n_4939));
OR2X1 g45454(.A (n_9717), .B (n_9666), .Y (n_11893));
CLKBUFX1 g45417(.A (n_11777), .Y (n_11762));
AOI22X1 g37815(.A0 (n_2558), .A1 (n_6380), .B0 (n_6664), .B1(n_2534), .Y (n_2527));
OAI21X1 g45459(.A0 (n_11908), .A1 (n_11914), .B0 (n_10481), .Y(n_11919));
NOR2X1 g40128(.A (n_2470), .B (n_2686), .Y (n_2107));
NOR2X1 g40129(.A (n_2477), .B (n_2801), .Y (n_2106));
NOR2X1 g45458(.A (n_11504), .B (dma_ack_i_b8_b), .Y (n_11907));
NOR2X1 g40120(.A (n_2470), .B (n_2831), .Y (n_2113));
NOR2X1 g40121(.A (n_2477), .B (n_2755), .Y (n_2111));
NOR2X1 g40122(.A (n_2477), .B (n_2786), .Y (n_2110));
NOR2X1 g40123(.A (n_1016), .B (n_2755), .Y (n_2757));
NOR2X1 g40124(.A (n_2470), .B (n_2794), .Y (n_2109));
NOR2X1 g40125(.A (n_2006), .B (n_2707), .Y (n_2114));
NOR2X1 g40126(.A (n_2189), .B (n_2720), .Y (n_2234));
NOR2X1 g40127(.A (n_2071), .B (n_2748), .Y (n_2108));
AOI21X1 g38447(.A0 (u6_mem_b3_b_147 ), .A1 (n_5100), .B0 (n_3350), .Y(n_4920));
MX2X1 g33129(.A (n_4713), .B (wb_din_662), .S0 (n_8611), .Y (n_8588));
MX2X1 g38633(.A (u4_mem_b0_b_121 ), .B (wb_din_691), .S0 (n_3765), .Y(n_3759));
AOI21X1 g45801(.A0 (n_12516), .A1 (n_12517), .B0 (n_12604), .Y(n_12520));
BUFX3 g40757(.A (n_938), .Y (n_4540));
NAND2X1 g45802(.A (n_6091), .B (n_12681), .Y (n_12516));
INVX4 g41531(.A (n_1320), .Y (n_3252));
INVX1 g41532(.A (n_1084), .Y (n_1320));
CLKBUFX3 g41533(.A (n_1084), .Y (n_2491));
INVX2 g41534(.A (n_532), .Y (n_1084));
NAND2X1 g41535(.A (n_12332), .B (n_12330), .Y (n_532));
NAND2X1 g41537(.A (u11_rp_b1_b ), .B (n_853), .Y (n_1121));
NAND2X1 g39009(.A (n_12839), .B (u4_mem_b0_b_107 ), .Y (n_3517));
NAND2X1 g39008(.A (u6_mem_b1_b_76 ), .B (n_12169), .Y (n_4249));
INVX4 g40755(.A (n_12752), .Y (n_1432));
NAND2X1 g39007(.A (n_12826), .B (u3_mem_b0_b_100 ), .Y (n_11719));
NAND2X1 g39006(.A (n_12369), .B (u6_mem_b0_b_120 ), .Y (n_3519));
NAND2X1 g41079(.A (n_697), .B (u26_ps_cnt_b0_b ), .Y (n_818));
NOR2X1 g39005(.A (n_3453), .B (n_2829), .Y (n_3520));
AOI22X1 g37809(.A0 (n_1756), .A1 (n_1628), .B0 (n_1627), .B1(n_1575), .Y (n_1629));
AOI22X1 g37808(.A0 (n_2558), .A1 (n_6331), .B0 (n_6565), .B1(n_1316), .Y (n_1317));
NAND2X1 g34502(.A (u5_mem_b1_b_79 ), .B (n_7870), .Y (n_7927));
OR2X1 g41522(.A (n_498), .B (n_459), .Y (n_976));
INVX1 g41521(.A (n_976), .Y (n_1122));
AOI22X1 g37801(.A0 (n_1756), .A1 (n_6388), .B0 (n_6500), .B1(n_1643), .Y (n_1638));
AOI22X1 g37800(.A0 (n_2502), .A1 (n_6398), .B0 (n_6654), .B1(n_1859), .Y (n_1639));
NAND2X1 g37803(.A (n_4183), .B (n_2700), .Y (n_5212));
AOI22X1 g37802(.A0 (n_6454), .A1 (n_1575), .B0 (n_6413), .B1(n_1831), .Y (n_1637));
AOI22X1 g37805(.A0 (n_1756), .A1 (n_1634), .B0 (n_1633), .B1(n_1643), .Y (n_1635));
MX2X1 g38749(.A (u3_mem_b0_b_115 ), .B (wb_din_685), .S0 (n_3807), .Y(n_3588));
AOI22X1 g37807(.A0 (n_81), .A1 (n_1575), .B0 (n_5494), .B1 (n_1831),.Y (n_1631));
NAND2X1 g37806(.A (n_3544), .B (n_2258), .Y (n_4581));
MX2X1 g33139(.A (wb_din_671), .B (oc1_cfg_976), .S0 (n_8538), .Y(n_8569));
MX2X1 g33138(.A (wb_din_670), .B (oc1_cfg_975), .S0 (n_8538), .Y(n_8570));
MX2X1 g38748(.A (u8_mem_b0_b_116 ), .B (wb_din_686), .S0 (n_3826), .Y(n_3589));
NAND2X1 g39001(.A (n_12825), .B (u3_mem_b0_b_111 ), .Y (n_3524));
NAND2X1 g39451(.A (n_3252), .B (u7_mem_b0_b_98 ), .Y (n_3171));
MX2X1 g33131(.A (n_4708), .B (wb_din_664), .S0 (n_8611), .Y (n_8584));
MX2X1 g33130(.A (n_4710), .B (wb_din_663), .S0 (n_8611), .Y (n_8586));
MX2X1 g33133(.A (n_4699), .B (wb_din_666), .S0 (n_8611), .Y (n_8579));
MX2X1 g33132(.A (n_4703), .B (wb_din_665), .S0 (n_8611), .Y (n_8581));
MX2X1 g33135(.A (n_11600), .B (wb_din_668), .S0 (n_8611), .Y(n_8575));
MX2X1 g33134(.A (ic0_cfg_1030), .B (wb_din_667), .S0 (n_8611), .Y(n_8577));
MX2X1 g33137(.A (wb_din), .B (n_862), .S0 (n_8538), .Y (n_8571));
MX2X1 g33136(.A (ic1_cfg_1034), .B (wb_din_669), .S0 (n_8611), .Y(n_8573));
MX2X1 g31151(.A (n_6897), .B (n_6895), .S0 (n_10277), .Y (n_10243));
MX2X1 g31150(.A (n_6022), .B (n_6021), .S0 (n_10315), .Y (n_10244));
MX2X1 g31153(.A (n_6887), .B (n_6886), .S0 (n_10308), .Y (n_10241));
MX2X1 g31152(.A (n_6914), .B (n_6912), .S0 (n_10308), .Y (n_10242));
MX2X1 g31155(.A (n_6019), .B (n_6018), .S0 (n_10565), .Y (n_10600));
MX2X1 g31154(.A (n_6910), .B (n_6909), .S0 (n_10250), .Y (n_10239));
MX2X1 g31157(.A (n_6907), .B (n_6905), .S0 (n_10235), .Y (n_10236));
MX2X1 g31156(.A (n_6561), .B (n_6559), .S0 (n_10235), .Y (n_10238));
MX2X1 g31159(.A (n_6603), .B (n_6601), .S0 (n_10137), .Y (n_10233));
MX2X1 g31158(.A (n_6006), .B (n_6005), .S0 (n_10137), .Y (n_10234));
OAI21X1 g30940(.A0 (n_1379), .A1 (o3_status), .B0 (n_9556), .Y(n_9584));
NAND2X1 g38878(.A (u8_mem_b3_b_140 ), .B (n_2468), .Y (n_2433));
MX2X1 g38743(.A (u8_mem_b0_b_108 ), .B (wb_din_678), .S0 (n_3826), .Y(n_3596));
OAI21X1 g30943(.A0 (n_1384), .A1 (o7_status), .B0 (n_9604), .Y(n_9643));
NAND2X1 g39457(.A (u6_mem_b1_b_67 ), .B (n_4253), .Y (n_11718));
AOI21X1 g38037(.A0 (u3_mem_b2_b_30 ), .A1 (n_4519), .B0 (n_2130), .Y(n_4518));
NAND2X1 g39849(.A (n_12826), .B (u3_mem_b0_b_98 ), .Y (n_2924));
AOI21X1 g38036(.A0 (u3_mem_b2_b_57 ), .A1 (n_4519), .B0 (n_2263), .Y(n_4520));
OAI21X1 g35898(.A0 (n_6085), .A1 (n_7187), .B0 (n_6785), .Y (n_7186));
OAI21X1 g35899(.A0 (n_6069), .A1 (n_7187), .B0 (n_5842), .Y (n_7184));
INVX1 g41109(.A (n_3522), .Y (n_1907));
OAI21X1 g35894(.A0 (n_5551), .A1 (n_7187), .B0 (n_5848), .Y (n_7016));
OAI21X1 g35896(.A0 (n_5549), .A1 (n_7187), .B0 (n_6817), .Y (n_7188));
OAI21X1 g35897(.A0 (n_5704), .A1 (n_7187), .B0 (n_5846), .Y (n_7093));
OAI21X1 g35890(.A0 (n_6075), .A1 (n_7187), .B0 (n_5854), .Y (n_7192));
OAI21X1 g35891(.A0 (n_6076), .A1 (n_7187), .B0 (n_6787), .Y (n_7190));
OAI21X1 g35892(.A0 (n_5552), .A1 (n_7187), .B0 (n_5852), .Y (n_6918));
OAI21X1 g35893(.A0 (n_6074), .A1 (n_7187), .B0 (n_5850), .Y (n_7189));
AOI21X1 g38033(.A0 (u3_mem_b2_b_54 ), .A1 (n_4519), .B0 (n_1971), .Y(n_4522));
NOR2X1 g39976(.A (n_867), .B (n_2748), .Y (n_2225));
MX2X1 g38744(.A (u3_mem_b0_b_110 ), .B (wb_din_680), .S0 (n_3807), .Y(n_3595));
XOR2X1 g37203(.A (n_1421), .B (n_4797), .Y (n_12838));
AOI21X1 g38254(.A0 (u8_mem_b1_b_60 ), .A1 (n_4387), .B0 (n_1981), .Y(n_4385));
OAI21X1 g36692(.A0 (n_5210), .A1 (n_5202), .B0 (n_6118), .Y (n_6096));
NAND2X1 g37753(.A (n_3087), .B (n_3224), .Y (n_4592));
INVX2 g35096(.A (n_7408), .Y (n_9307));
INVX1 g35097(.A (n_7408), .Y (n_9288));
INVX1 g35090(.A (n_7408), .Y (n_9202));
INVX1 g35092(.A (n_7408), .Y (n_9230));
INVX1 g35093(.A (n_7408), .Y (n_9205));
MX2X1 g37207(.A (u9_mem_b1_b_140 ), .B (n_4776), .S0 (n_4783), .Y(n_4794));
XOR2X1 g37206(.A (u8_wp_b0_b ), .B (n_3992), .Y (n_3993));
NAND2X1 g37757(.A (n_3274), .B (n_2982), .Y (n_4591));
AOI22X1 g37756(.A0 (n_2558), .A1 (n_2539), .B0 (n_2538), .B1 (n_940),.Y (n_2540));
NAND2X1 g38929(.A (u7_mem_b3_b_144 ), .B (n_1546), .Y (n_1527));
NAND2X1 g38928(.A (u7_mem_b3_b_128 ), .B (n_1538), .Y (n_1528));
AND2X1 g35270(.A (n_4846), .B (u2_sync_resume), .Y (n_5628));
NOR2X1 g35271(.A (n_7141), .B (n_11762), .Y (n_7371));
NAND2X1 g35272(.A (n_6674), .B (n_7331), .Y (n_7488));
NAND2X1 g35273(.A (n_6678), .B (n_7330), .Y (n_7487));
NAND2X1 g35274(.A (n_6699), .B (n_7336), .Y (n_7486));
NOR2X1 g35275(.A (n_7143), .B (n_11563), .Y (n_7369));
NAND2X1 g35276(.A (n_7112), .B (n_7335), .Y (n_7485));
NAND2X1 g35277(.A (n_6685), .B (n_7333), .Y (n_7484));
NAND2X1 g35278(.A (n_6690), .B (n_7332), .Y (n_7483));
NAND2X1 g35279(.A (n_7329), .B (n_6697), .Y (n_7482));
NAND2X1 g40724(.A (n_8536), .B (n_571), .Y (n_9645));
CLKBUFX1 g40725(.A (n_940), .Y (n_1839));
NAND2X1 g40722(.A (n_706), .B (u6_wp_b1_b ), .Y (n_941));
NOR2X1 g40723(.A (n_8536), .B (n_571), .Y (n_9766));
INVX1 g40720(.A (n_1176), .Y (n_2144));
NAND2X1 g39859(.A (n_12721), .B (u3_mem_b0_b_92 ), .Y (n_2917));
OAI21X1 g33041(.A0 (n_7247), .A1 (n_7087), .B0 (n_12504), .Y(n_10204));
INVX1 g42387(.A (n_9833), .Y (n_10921));
INVX1 g39857(.A (n_4753), .Y (n_2918));
INVX1 g43038(.A (n_1873), .Y (n_1870));
CLKBUFX1 g43031(.A (n_1873), .Y (n_1875));
NAND2X1 g39851(.A (n_4560), .B (in_slt_444), .Y (n_2922));
NAND2X1 g39852(.A (n_11789), .B (u8_mem_b0_b_92 ), .Y (n_12844));
NAND3X1 g39151(.A (u8_mem_b0_b_106 ), .B (n_12280), .C (n_691), .Y(n_1493));
NAND2X1 g39150(.A (u7_mem_b1_b_87 ), .B (n_4225), .Y (n_4223));
INVX4 g39157(.A (n_1453), .Y (n_6972));
NAND2X1 g38871(.A (u8_mem_b3_b_122 ), .B (n_2468), .Y (n_2435));
AOI22X1 g40415(.A0 (u13_intm_r_b5_b ), .A1 (u13_ints_r_b5_b ), .B0(u13_intm_r_b6_b ), .B1 (u13_ints_r_b6_b ), .Y (n_728));
MX2X1 g34059(.A (u6_mem_b0_b_110 ), .B (n_3609), .S0 (n_7505), .Y(n_8770));
MX2X1 g34058(.A (u6_mem_b0_b_91 ), .B (n_3630), .S0 (n_7505), .Y(n_8772));
MX2X1 g34057(.A (u6_mem_b0_b_109 ), .B (n_3573), .S0 (n_7505), .Y(n_9411));
MX2X1 g34056(.A (u6_mem_b0_b_108 ), .B (n_3674), .S0 (n_7505), .Y(n_8773));
MX2X1 g34055(.A (u6_mem_b0_b_107 ), .B (n_3576), .S0 (n_7505), .Y(n_8775));
MX2X1 g34054(.A (u6_mem_b0_b_106 ), .B (n_3675), .S0 (n_7505), .Y(n_9412));
MX2X1 g34053(.A (u6_mem_b0_b_105 ), .B (n_3676), .S0 (n_7505), .Y(n_8776));
MX2X1 g34052(.A (u6_mem_b0_b_104 ), .B (n_3567), .S0 (n_7505), .Y(n_9413));
MX2X1 g34051(.A (u6_mem_b0_b_103 ), .B (n_3679), .S0 (n_7505), .Y(n_9414));
MX2X1 g34050(.A (u6_mem_b0_b_102 ), .B (n_3681), .S0 (n_7505), .Y(n_8778));
INVX1 g41858(.A (u10_mem_b0_b_158 ), .Y (n_5962));
AOI21X1 g45525(.A0 (n_12131), .A1 (n_12132), .B0 (n_12145), .Y(n_12135));
INVX4 g40596(.A (wb_din_668), .Y (n_2772));
NAND2X1 g29929(.A (n_11158), .B (u16_u3_dma_req_r1), .Y (n_11182));
NAND2X1 g29928(.A (n_11124), .B (u16_u2_dma_req_r1), .Y (n_11172));
NAND2X1 g29927(.A (n_11159), .B (u16_u1_dma_req_r1), .Y (n_11183));
NAND2X1 g29926(.A (n_11125), .B (u16_u0_dma_req_r1), .Y (n_11173));
AOI21X1 g38350(.A0 (u5_mem_b3_b_122 ), .A1 (n_4996), .B0 (n_2975), .Y(n_4987));
AOI21X1 g38351(.A0 (u5_mem_b3_b_141 ), .A1 (n_5000), .B0 (n_3449), .Y(n_4986));
AOI21X1 g38352(.A0 (u5_mem_b3_b_142 ), .A1 (n_5000), .B0 (n_3053), .Y(n_4985));
AOI21X1 g38353(.A0 (u5_mem_b3_b_143 ), .A1 (n_4996), .B0 (n_3131), .Y(n_4984));
AOI21X1 g38354(.A0 (u5_mem_b3_b_144 ), .A1 (n_4996), .B0 (n_3129), .Y(n_4983));
AOI21X1 g38356(.A0 (u5_mem_b3_b_146 ), .A1 (n_4996), .B0 (n_3001), .Y(n_4981));
AOI21X1 g38357(.A0 (u5_mem_b3_b_147 ), .A1 (n_4996), .B0 (n_3006), .Y(n_4980));
INVX1 g37126(.A (n_6783), .Y (n_6069));
NAND4X1 g37127(.A (n_11514), .B (n_3142), .C (n_11515), .D (n_2414),.Y (n_6783));
NOR2X1 g37124(.A (n_5413), .B (n_6649), .Y (n_4804));
NOR2X1 g37125(.A (n_5410), .B (n_6649), .Y (n_4803));
NAND4X1 g37122(.A (n_3135), .B (n_2917), .C (n_3405), .D (n_1378), .Y(n_6184));
MX2X1 g38603(.A (u3_mem_b0_b ), .B (wb_din), .S0 (n_3807), .Y(n_3808));
NAND4X1 g37120(.A (n_3355), .B (n_2861), .C (n_2295), .D (n_2381), .Y(n_5893));
INVX1 g37121(.A (n_6184), .Y (n_5668));
OAI21X1 g33728(.A0 (n_4936), .A1 (n_9182), .B0 (n_7801), .Y (n_9158));
OAI21X1 g33729(.A0 (n_4935), .A1 (n_9077), .B0 (n_7800), .Y (n_9157));
NAND2X1 g38877(.A (u5_mem_b3_b_134 ), .B (n_1543), .Y (n_1534));
OAI21X1 g33724(.A0 (n_4939), .A1 (n_9165), .B0 (n_7806), .Y (n_9166));
OAI21X1 g33725(.A0 (n_5054), .A1 (n_9087), .B0 (n_7804), .Y (n_9164));
OAI21X1 g33726(.A0 (n_4937), .A1 (n_9161), .B0 (n_7803), .Y (n_9162));
OAI21X1 g33727(.A0 (n_5140), .A1 (n_9110), .B0 (n_7802), .Y (n_9160));
OAI21X1 g33720(.A0 (n_4940), .A1 (n_9170), .B0 (n_7810), .Y (n_9171));
OAI21X1 g33721(.A0 (n_5008), .A1 (n_9165), .B0 (n_7809), .Y (n_9169));
OAI21X1 g33722(.A0 (n_5011), .A1 (n_9139), .B0 (n_7808), .Y (n_9168));
OAI21X1 g33723(.A0 (n_5020), .A1 (n_9087), .B0 (n_7807), .Y (n_9167));
NAND2X1 g38876(.A (u7_mem_b3_b_148 ), .B (n_1546), .Y (n_1535));
INVX1 g42812(.A (n_454), .Y (n_4701));
INVX1 g42810(.A (u10_mem_b2_b_117 ), .Y (n_2542));
INVX1 g42811(.A (u11_mem_b0_b_178 ), .Y (n_1592));
NAND2X1 g36529(.A (n_12111), .B (n_12115), .Y (n_6220));
NAND2X1 g36528(.A (n_6153), .B (n_6259), .Y (n_6221));
NOR2X1 g36525(.A (o6_status), .B (n_2485), .Y (n_5438));
NAND2X1 g36524(.A (n_2566), .B (n_4834), .Y (n_5964));
NAND2X1 g36527(.A (n_5829), .B (n_784), .Y (n_5830));
NAND2X1 g36526(.A (n_1772), .B (n_4080), .Y (n_5636));
NAND2X1 g36521(.A (n_6816), .B (n_5833), .Y (n_5834));
NAND2X1 g36520(.A (n_6781), .B (n_784), .Y (n_6782));
NAND2X1 g36523(.A (n_6779), .B (n_6816), .Y (n_6780));
MX2X1 g31095(.A (n_6029), .B (n_6028), .S0 (n_10450), .Y (n_10652));
INVX2 g42978(.A (n_1481), .Y (n_11144));
INVX1 g42603(.A (u3_rp_b2_b ), .Y (n_601));
INVX1 g42602(.A (n_601), .Y (n_763));
INVX1 g42977(.A (u9_mem_b3_b_71 ), .Y (n_6581));
INVX1 g42976(.A (u10_mem_b0_b_150 ), .Y (n_5949));
INVX1 g42970(.A (u9_mem_b3_b_82 ), .Y (n_5369));
INVX1 g42605(.A (u9_mem_b1_b_139 ), .Y (n_1679));
INVX1 g42604(.A (u3_rp_b2_b ), .Y (n_63));
NAND2X1 g41778(.A (u9_rp_b1_b ), .B (u9_wp_b2_b ), .Y (n_984));
INVX4 g40638(.A (wb_din_683), .Y (n_2684));
OR2X1 g41776(.A (n_1355), .B (n_5827), .Y (n_1356));
AND2X1 g41777(.A (n_671), .B (n_924), .Y (n_9614));
OR2X1 g41775(.A (n_1100), .B (n_5825), .Y (n_1101));
AOI22X1 g36749(.A0 (n_5630), .A1 (u2_to_cnt_b1_b ), .B0 (n_5629), .B1(n_795), .Y (n_5404));
XOR2X1 g36748(.A (n_1188), .B (n_1160), .Y (n_2611));
INVX1 g41850(.A (u10_mem_b0_b_175 ), .Y (n_1677));
MX2X1 g36740(.A (u10_mem_b1_b_136 ), .B (n_5418), .S0 (n_5407), .Y(n_5408));
XOR2X1 g36743(.A (u26_cnt_b2_b ), .B (n_793), .Y (n_1821));
MX2X1 g36742(.A (u11_mem_b1_b_137 ), .B (n_5410), .S0 (n_5405), .Y(n_5406));
XOR2X1 g36745(.A (u2_res_cnt_b2_b ), .B (n_1277), .Y (n_1818));
XOR2X1 g36744(.A (n_1819), .B (n_1553), .Y (n_1820));
XOR2X1 g36747(.A (n_786), .B (n_1164), .Y (n_2612));
XOR2X1 g36746(.A (n_1157), .B (n_1438), .Y (n_4072));
INVX1 g36999(.A (n_6224), .Y (n_5703));
OAI21X1 g30966(.A0 (n_4754), .A1 (n_10747), .B0 (n_9995), .Y(n_10748));
OAI21X1 g30965(.A0 (n_4789), .A1 (n_10747), .B0 (n_10059), .Y(n_10750));
OAI21X1 g30964(.A0 (n_4794), .A1 (n_10738), .B0 (n_10060), .Y(n_10751));
OAI21X1 g30963(.A0 (n_5342), .A1 (n_10450), .B0 (n_10058), .Y(n_10752));
OAI21X1 g30962(.A0 (n_4790), .A1 (n_10738), .B0 (n_10062), .Y(n_10753));
OAI21X1 g30961(.A0 (n_4791), .A1 (n_10747), .B0 (n_10063), .Y(n_10754));
OAI21X1 g30960(.A0 (n_5731), .A1 (n_10747), .B0 (n_9991), .Y(n_10755));
NAND2X1 g39438(.A (u3_mem_b1_b_70 ), .B (n_12753), .Y (n_11722));
NAND2X1 g39439(.A (u3_mem_b1_b_60 ), .B (n_3316), .Y (n_3183));
OAI21X1 g30969(.A0 (n_4786), .A1 (n_10747), .B0 (n_10055), .Y(n_10743));
OAI21X1 g30968(.A0 (n_4750), .A1 (n_10738), .B0 (n_10056), .Y(n_10744));
OAI21X1 g33922(.A0 (n_4400), .A1 (n_8891), .B0 (n_7601), .Y (n_8918));
NAND2X1 g34603(.A (u6_mem_b1_b_73 ), .B (n_7758), .Y (n_7825));
NAND2X1 g34600(.A (u6_mem_b1_b_70 ), .B (n_7758), .Y (n_7830));
NAND2X1 g34601(.A (u6_mem_b1_b_71 ), .B (n_7758), .Y (n_7828));
NAND2X1 g34606(.A (u6_mem_b1_b_76 ), .B (n_7758), .Y (n_7822));
NAND2X1 g34607(.A (u6_mem_b1_b_77 ), .B (n_7758), .Y (n_7821));
NAND2X1 g34604(.A (u6_mem_b1_b_74 ), .B (n_7758), .Y (n_7824));
NAND2X1 g34605(.A (u6_mem_b1_b_75 ), .B (n_7758), .Y (n_7823));
NAND2X1 g34608(.A (u6_mem_b1_b_78 ), .B (n_7758), .Y (n_7819));
NAND2X1 g34609(.A (u3_mem_b1_b_65 ), .B (n_8101), .Y (n_7818));
MX2X1 g31217(.A (n_6438), .B (n_6437), .S0 (n_10513), .Y (n_10494));
MX2X1 g31214(.A (n_6449), .B (n_6448), .S0 (n_10513), .Y (n_10508));
MX2X1 g31215(.A (n_6446), .B (n_6445), .S0 (n_10513), .Y (n_10501));
MX2X1 g31212(.A (n_5973), .B (n_501), .S0 (n_10315), .Y (n_10190));
MX2X1 g31213(.A (n_5971), .B (n_406), .S0 (n_10315), .Y (n_10187));
MX2X1 g31210(.A (n_6452), .B (n_502), .S0 (n_10315), .Y (n_10197));
MX2X1 g31211(.A (n_5975), .B (n_5974), .S0 (n_10315), .Y (n_10194));
MX2X1 g31218(.A (n_6435), .B (n_6434), .S0 (n_10513), .Y (n_10489));
MX2X1 g31219(.A (n_6531), .B (n_6530), .S0 (n_10839), .Y (n_10838));
AOI22X1 g40410(.A0 (u13_intm_r_b14_b ), .A1 (u13_ints_r_b14_b ), .B0(u13_intm_r_b16_b ), .B1 (u13_ints_r_b16_b ), .Y (n_732));
NAND2X1 g39388(.A (u5_mem_b1_b_75 ), .B (n_3257), .Y (n_3218));
NAND2X1 g39389(.A (n_3259), .B (u5_mem_b0_b_106 ), .Y (n_11966));
INVX1 g42473(.A (u10_mem_b2_b_104 ), .Y (n_6030));
NOR2X1 g39384(.A (n_1484), .B (n_760), .Y (n_1485));
NOR2X1 g39385(.A (n_713), .B (u26_cnt_b0_b ), .Y (n_1777));
NAND2X1 g39386(.A (u4_mem_b2_b_30 ), .B (n_12079), .Y (n_2314));
NOR2X1 g39387(.A (n_3332), .B (n_2763), .Y (n_3220));
NAND2X1 g39380(.A (in_slt_411), .B (n_3415), .Y (n_3223));
NAND2X1 g39381(.A (u5_mem_b1_b_74 ), .B (n_3236), .Y (n_12842));
NAND2X1 g39383(.A (u5_mem_b2_b_43 ), .B (n_12823), .Y (n_12041));
BUFX3 g40771(.A (n_945), .Y (n_4519));
BUFX3 g45579(.A (n_12364), .Y (n_12204));
OAI21X1 g33948(.A0 (n_4494), .A1 (n_8438), .B0 (n_7579), .Y (n_8881));
OAI21X1 g33519(.A0 (n_4460), .A1 (n_9326), .B0 (n_8039), .Y (n_8328));
NAND2X1 g34669(.A (u6_mem_b3_b_134 ), .B (n_7758), .Y (n_7755));
NAND2X1 g34237(.A (u3_mem_b1_b_61 ), .B (n_8101), .Y (n_8169));
AOI22X1 g35710(.A0 (n_6686), .A1 (i6_dout_641), .B0 (i4_dout_610),.B1 (n_7297), .Y (n_6674));
INVX4 g41363(.A (n_1851), .Y (n_6341));
NAND2X1 g34236(.A (u8_mem_b2_b_35 ), .B (n_7976), .Y (n_8171));
OAI21X1 g33515(.A0 (n_4464), .A1 (n_8333), .B0 (n_8045), .Y (n_8334));
CLKBUFX1 g35240(.A (o9_we), .Y (n_7396));
OAI21X1 g33514(.A0 (n_4475), .A1 (n_8333), .B0 (n_8046), .Y (n_8336));
BUFX3 g41584(.A (n_5059), .Y (n_5100));
INVX4 g45893(.A (n_12621), .Y (n_12622));
NAND2X1 g34660(.A (u6_mem_b2_b_33 ), .B (n_7758), .Y (n_7765));
INVX4 g45890(.A (n_1429), .Y (n_12619));
INVX2 g40631(.A (wb_din_677), .Y (n_2735));
NAND2X1 g45896(.A (n_12369), .B (u6_mem_b0_b_104 ), .Y (n_12624));
NOR2X1 g45895(.A (n_11579), .B (n_192), .Y (n_12620));
NAND2X1 g34661(.A (u6_mem_b2_b_34 ), .B (n_7758), .Y (n_7764));
NAND3X1 g45899(.A (n_12627), .B (n_12636), .C (u7_rp_b0_b ), .Y(n_12630));
NAND2X1 g45898(.A (n_12630), .B (n_12631), .Y (n_12632));
NAND2X1 g34662(.A (u6_mem_b2_b_35 ), .B (n_7758), .Y (n_7763));
NAND2X1 g34663(.A (u6_mem_b2_b_36 ), .B (n_7758), .Y (n_7762));
AOI21X1 g30030(.A0 (n_9551), .A1 (n_9695), .B0 (n_10087), .Y(n_10406));
OAI21X1 g33944(.A0 (n_4331), .A1 (n_8433), .B0 (n_7805), .Y (n_8886));
OAI21X1 g33945(.A0 (n_4344), .A1 (n_8464), .B0 (n_7582), .Y (n_8885));
NAND2X1 g34666(.A (u6_mem_b3_b_131 ), .B (n_7758), .Y (n_7759));
NAND2X1 g34667(.A (u6_mem_b3_b_132 ), .B (n_7758), .Y (n_7757));
BUFX3 g40711(.A (n_941), .Y (n_4504));
INVX4 g40815(.A (n_877), .Y (n_1859));
AOI21X1 g38167(.A0 (u4_mem_b2_b_56 ), .A1 (n_4439), .B0 (n_2012), .Y(n_4420));
AOI21X1 g38166(.A0 (u4_mem_b2_b_55 ), .A1 (n_4439), .B0 (n_1970), .Y(n_4421));
AOI21X1 g38165(.A0 (u7_mem_b1_b_74 ), .A1 (n_5118), .B0 (n_2670), .Y(n_5110));
AOI21X1 g38164(.A0 (u4_mem_b2_b_54 ), .A1 (n_4439), .B0 (n_2048), .Y(n_4422));
AOI21X1 g38163(.A0 (u4_mem_b2_b_53 ), .A1 (n_4439), .B0 (n_2484), .Y(n_4423));
AOI21X1 g38162(.A0 (u7_mem_b2_b_40 ), .A1 (n_4509), .B0 (n_1994), .Y(n_4424));
AOI21X1 g38161(.A0 (u4_mem_b2_b_52 ), .A1 (n_4439), .B0 (n_1998), .Y(n_4425));
AOI21X1 g38160(.A0 (u4_mem_b2_b_51 ), .A1 (n_4439), .B0 (n_2100), .Y(n_4426));
NAND2X1 g39232(.A (in_slt_410), .B (n_3415), .Y (n_3348));
NAND2X1 g39950(.A (u8_mem_b2_b_40 ), .B (n_2366), .Y (n_11454));
AOI21X1 g38169(.A0 (u4_mem_b2_b_57 ), .A1 (n_4439), .B0 (n_2024), .Y(n_4419));
AOI21X1 g38168(.A0 (u6_mem_b3_b_124 ), .A1 (n_5100), .B0 (n_3507), .Y(n_5109));
INVX1 g40777(.A (n_1172), .Y (n_2085));
NAND2X1 g36408(.A (n_7049), .B (n_7048), .Y (n_6268));
NAND2X1 g36409(.A (n_6842), .B (n_6841), .Y (n_5902));
NOR2X1 g40142(.A (n_867), .B (n_2720), .Y (n_2226));
NAND2X1 g36406(.A (n_5859), .B (n_3559), .Y (n_5904));
NOR2X1 g40140(.A (n_935), .B (n_2712), .Y (n_2095));
NOR2X1 g40141(.A (n_2093), .B (n_2794), .Y (n_2094));
NOR2X1 g40146(.A (n_2477), .B (n_2831), .Y (n_2484));
NOR2X1 g40147(.A (n_2801), .B (n_2067), .Y (n_2091));
NOR2X1 g40144(.A (n_2751), .B (n_2716), .Y (n_2752));
NAND2X1 g36407(.A (n_6836), .B (u8_wp_b1_b ), .Y (n_5903));
NOR2X1 g40149(.A (n_1082), .B (n_2744), .Y (n_2746));
AOI21X1 g38291(.A0 (u5_mem_b1_b_61 ), .A1 (n_5037), .B0 (n_2672), .Y(n_5021));
AOI21X1 g38290(.A0 (u5_mem_b1_b_88 ), .A1 (n_5048), .B0 (n_2806), .Y(n_5022));
AOI21X1 g38293(.A0 (u5_mem_b1_b_89 ), .A1 (n_5037), .B0 (n_2828), .Y(n_5018));
AOI21X1 g38292(.A0 (u6_mem_b1_b_86 ), .A1 (n_5019), .B0 (n_2764), .Y(n_5020));
AOI21X1 g38295(.A0 (u5_mem_b1_b_62 ), .A1 (n_5037), .B0 (n_2800), .Y(n_5016));
AOI21X1 g38294(.A0 (u5_mem_b1_b_90 ), .A1 (n_5037), .B0 (n_2719), .Y(n_5017));
AOI21X1 g38297(.A0 (u5_mem_b1_b_64 ), .A1 (n_5037), .B0 (n_2746), .Y(n_5014));
AOI21X1 g38296(.A0 (u5_mem_b1_b_63 ), .A1 (n_5037), .B0 (n_2967), .Y(n_5015));
AOI21X1 g38299(.A0 (u5_mem_b1_b_66 ), .A1 (n_5037), .B0 (n_2835), .Y(n_5012));
NAND2X1 g31685(.A (n_1591), .B (n_10376), .Y (n_10377));
INVX1 g42374(.A (u10_wp_b1_b ), .Y (n_708));
INVX4 g45432(.A (n_11797), .Y (n_11798));
INVX1 g41927(.A (ic0_int_set_720), .Y (n_739));
NAND2X1 g37970(.A (n_2915), .B (n_2935), .Y (n_5173));
NAND2X1 g34444(.A (u4_mem_b3_b_141 ), .B (n_7984), .Y (n_7970));
AOI22X1 g34917(.A0 (n_5630), .A1 (u2_to_cnt_b3_b ), .B0 (n_5629), .B1(n_4100), .Y (n_5631));
NAND2X1 g37975(.A (n_2409), .B (n_2870), .Y (n_5170));
OAI21X1 g33635(.A0 (n_5010), .A1 (n_9286), .B0 (n_7907), .Y (n_9275));
OAI21X1 g33490(.A0 (n_5066), .A1 (n_8383), .B0 (n_8081), .Y (n_8363));
AOI22X1 g37355(.A0 (n_4729), .A1 (oc4_cfg_1010), .B0 (n_5591), .B1(ic0_cfg_1030), .Y (n_4698));
AOI22X1 g37354(.A0 (n_5272), .A1 (u13_intm_r_b7_b ), .B0 (n_5277), .B1(crac_din_698), .Y (n_5260));
AOI22X1 g37357(.A0 (n_4729), .A1 (n_8182), .B0 (n_5591), .B1(n_11600), .Y (n_4697));
OAI21X1 g33491(.A0 (n_5127), .A1 (n_8383), .B0 (n_8082), .Y (n_8362));
AOI22X1 g37351(.A0 (n_4729), .A1 (n_8188), .B0 (n_5591), .B1(n_4703), .Y (n_4704));
AOI22X1 g37350(.A0 (n_5272), .A1 (u13_intm_r_b5_b ), .B0 (n_5277), .B1(crac_din_696), .Y (n_5263));
AOI22X1 g37352(.A0 (n_5272), .A1 (u13_intm_r_b6_b ), .B0 (n_5277), .B1(crac_din_697), .Y (n_5261));
AOI22X1 g37829(.A0 (n_6018), .A1 (n_2553), .B0 (n_6000), .B1(n_1316), .Y (n_2523));
AOI22X1 g37828(.A0 (n_122), .A1 (n_1575), .B0 (n_5522), .B1 (n_1831),.Y (n_1602));
AOI22X1 g37359(.A0 (n_4729), .A1 (oc5_cfg_1014), .B0 (n_5591), .B1(ic1_cfg_1034), .Y (n_4695));
AOI22X1 g37358(.A0 (n_5272), .A1 (u13_intm_r_b9_b ), .B0 (n_5277), .B1(crac_din_700), .Y (n_5256));
MX2X1 g33113(.A (n_11564), .B (wb_din), .S0 (n_8611), .Y (n_8624));
MX2X1 g33112(.A (crac_out_876), .B (wb_din_691), .S0 (n_8643), .Y(n_8626));
MX2X1 g33111(.A (crac_out_867), .B (wb_din_682), .S0 (n_8643), .Y(n_8627));
MX2X1 g33110(.A (crac_out_866), .B (wb_din_681), .S0 (n_8643), .Y(n_8628));
MX2X1 g33117(.A (n_4734), .B (wb_din_673), .S0 (n_8611), .Y (n_8616));
MX2X1 g33116(.A (n_4736), .B (wb_din_672), .S0 (n_8611), .Y (n_8618));
MX2X1 g33115(.A (n_4690), .B (wb_din_671), .S0 (n_8611), .Y (n_8620));
MX2X1 g33114(.A (n_4738), .B (wb_din_670), .S0 (n_8611), .Y (n_8622));
INVX4 g41549(.A (n_12621), .Y (n_2465));
MX2X1 g33119(.A (ic1_cfg_1040), .B (wb_din_675), .S0 (n_8611), .Y(n_8610));
OAI21X1 g36198(.A0 (n_6836), .A1 (u8_wp_b1_b ), .B0 (n_5903), .Y(n_6837));
ADDHX1 g36199(.A (n_686), .B (u10_wp_b2_b ), .CO (n_1559), .S(n_1560));
INVX1 g43029(.A (n_1875), .Y (n_11083));
XOR2X1 g36194(.A (n_657), .B (n_5942), .Y (n_5944));
OAI21X1 g36195(.A0 (n_7049), .A1 (n_7048), .B0 (n_6268), .Y (n_7050));
OAI21X1 g36196(.A0 (n_6842), .A1 (n_6841), .B0 (n_5902), .Y (n_6843));
OAI21X1 g36197(.A0 (n_6839), .A1 (n_6838), .B0 (n_5901), .Y (n_6840));
XOR2X1 g36190(.A (n_799), .B (n_1788), .Y (n_4841));
XOR2X1 g36191(.A (n_1418), .B (n_1267), .Y (n_4091));
XOR2X1 g36192(.A (n_1422), .B (n_1265), .Y (n_4090));
XOR2X1 g36193(.A (n_614), .B (n_6328), .Y (n_6330));
MX2X1 g31179(.A (n_6516), .B (n_6515), .S0 (n_10839), .Y (n_10844));
MX2X1 g31178(.A (n_6518), .B (n_6517), .S0 (n_10513), .Y (n_10561));
NAND2X1 g38912(.A (u4_mem_b3_b_127 ), .B (n_3546), .Y (n_3534));
MX2X1 g31173(.A (n_6564), .B (n_6562), .S0 (n_10137), .Y (n_10217));
MX2X1 g31172(.A (n_6567), .B (n_6565), .S0 (n_10137), .Y (n_10219));
MX2X1 g31171(.A (n_6571), .B (n_6569), .S0 (n_10137), .Y (n_10220));
MX2X1 g31170(.A (n_6574), .B (n_6572), .S0 (n_10137), .Y (n_10221));
MX2X1 g31177(.A (n_6520), .B (n_6519), .S0 (n_10513), .Y (n_10562));
MX2X1 g31176(.A (n_6523), .B (n_6522), .S0 (n_10513), .Y (n_10563));
MX2X1 g31175(.A (n_6001), .B (n_6000), .S0 (n_10565), .Y (n_10564));
MX2X1 g31174(.A (n_6004), .B (n_6002), .S0 (n_10137), .Y (n_10216));
MX2X1 g36088(.A (n_6495), .B (n_6539), .S0 (n_6898), .Y (n_6496));
NOR2X1 g40982(.A (n_1923), .B (n_1419), .Y (n_1420));
CLKBUFX3 g41110(.A (n_11851), .Y (n_3522));
NOR2X1 g39148(.A (n_3453), .B (n_3008), .Y (n_3417));
NOR2X1 g40983(.A (n_11585), .B (n_1417), .Y (n_1418));
NOR2X1 g40025(.A (n_945), .B (n_2729), .Y (n_2191));
NOR2X1 g40980(.A (n_1033), .B (n_798), .Y (n_799));
INVX1 g41926(.A (u10_mem_b2_b_102 ), .Y (n_6660));
AND2X1 g40981(.A (n_621), .B (wb_addr_i_b3_b), .Y (n_1225));
NAND2X1 g38910(.A (u5_mem_b3_b_137 ), .B (n_3543), .Y (n_2406));
NOR2X1 g40285(.A (n_2767), .B (n_1985), .Y (n_1989));
NOR2X1 g40284(.A (n_2689), .B (n_2755), .Y (n_2680));
INVX2 g35077(.A (n_7414), .Y (n_8318));
OR2X1 g32970_dup(.A (n_9719), .B (n_9668), .Y (n_11892));
NOR2X1 g40287(.A (n_2742), .B (n_2744), .Y (n_2679));
NOR2X1 g40286(.A (n_2755), .B (n_2118), .Y (n_1988));
INVX1 g45450(.A (n_11852), .Y (n_11853));
INVX4 g41116(.A (n_11852), .Y (n_4130));
NOR2X1 g40281(.A (n_1082), .B (n_2684), .Y (n_2685));
NOR2X1 g40280(.A (n_2154), .B (n_2864), .Y (n_1990));
NOR2X1 g35832(.A (n_7353), .B (n_5268), .Y (n_7111));
NAND2X1 g39144(.A (in_slt_410), .B (n_2368), .Y (n_4749));
AND2X1 g35833(.A (n_1285), .B (n_5248), .Y (n_5361));
INVX1 g42014(.A (u10_mem_b1_b_135 ), .Y (n_501));
NOR2X1 g40282(.A (n_1147), .B (n_2741), .Y (n_2683));
NOR2X1 g35830(.A (n_4830), .B (n_2622), .Y (n_5613));
NAND2X1 g38916(.A (u5_mem_b3_b_143 ), .B (n_3543), .Y (n_2404));
INVX1 g42011(.A (u9_mem_b0_b_157 ), .Y (n_6394));
NOR2X1 g35836(.A (n_4835), .B (n_2619), .Y (n_5612));
INVX1 g40748(.A (n_3316), .Y (n_1918));
NOR2X1 g35837(.A (n_4082), .B (n_2618), .Y (n_5383));
NAND2X1 g40708(.A (n_8565), .B (n_942), .Y (n_9647));
NOR2X1 g40709(.A (n_3559), .B (u5_rp_b3_b ), .Y (n_785));
NAND3X1 g35834(.A (n_4084), .B (n_731), .C (n_577), .Y (n_5444));
INVX8 g35212(.A (o9_we), .Y (n_7976));
INVX1 g40701(.A (n_1434), .Y (n_3334));
NAND2X1 g38917(.A (u6_mem_b3_b_142 ), .B (n_2465), .Y (n_2403));
CLKBUFX3 g40705(.A (n_1178), .Y (n_2366));
INVX2 g40706(.A (n_714), .Y (n_1178));
NAND2X2 g40707(.A (n_12274), .B (n_691), .Y (n_714));
INVX1 g41938(.A (n_8182), .Y (n_11033));
NAND2X1 g39173(.A (u8_mem_b1_b_81 ), .B (n_12291), .Y (n_3404));
NAND2X1 g39172(.A (u4_mem_b2_b_45 ), .B (n_12079), .Y (n_2350));
OR2X1 g39171(.A (n_12145), .B (n_6824), .Y (n_1460));
NAND2X1 g39170(.A (u3_mem_b2_b_30 ), .B (n_12619), .Y (n_3405));
NOR2X1 g39177(.A (n_3089), .B (n_2684), .Y (n_3400));
NAND2X1 g39176(.A (u4_mem_b2_b_58 ), .B (n_12079), .Y (n_3401));
NAND2X1 g39175(.A (u3_mem_b1_b ), .B (n_3316), .Y (n_12831));
NAND2X1 g39174(.A (u4_mem_b1_b_80 ), .B (n_12265), .Y (n_4219));
INVX1 g43051(.A (u10_mem_b3_b_61 ), .Y (n_6569));
INVX1 g43050(.A (u9_mem_b0_b_154 ), .Y (n_6852));
NAND2X1 g39179(.A (n_12839), .B (u4_mem_b0_b_120 ), .Y (n_2950));
NAND2X1 g39178(.A (u4_mem_b1_b_89 ), .B (n_12267), .Y (n_4218));
INVX1 g43055(.A (u10_mem_b3_b_78 ), .Y (n_5518));
INVX1 g43057(.A (u9_mem_b3_b_64 ), .Y (n_6559));
INVX1 g43056(.A (u10_mem_b2_b_94 ), .Y (n_6607));
NAND2X1 g38915(.A (u8_mem_b3_b_127 ), .B (n_2468), .Y (n_1881));
INVX1 g42232(.A (u11_mem_b3_b_87 ), .Y (n_5522));
NAND2X1 g38819(.A (u4_mem_b3_b_123 ), .B (n_4258), .Y (n_4257));
INVX1 g42589(.A (u9_mem_b3_b_84 ), .Y (n_5347));
INVX1 g41934(.A (n_8182), .Y (n_11025));
MX2X1 g34039(.A (u5_mem_b0_b_93 ), .B (n_3697), .S0 (n_7496), .Y(n_8786));
MX2X1 g34038(.A (u5_mem_b0_b_121 ), .B (n_3698), .S0 (n_7496), .Y(n_9421));
MX2X1 g34031(.A (u5_mem_b0_b_115 ), .B (n_3712), .S0 (n_7496), .Y(n_8794));
MX2X1 g34030(.A (u5_mem_b0_b_114 ), .B (n_3714), .S0 (n_7496), .Y(n_9422));
MX2X1 g34032(.A (u5_mem_b0_b_116 ), .B (n_3709), .S0 (n_7496), .Y(n_8793));
MX2X1 g34035(.A (u5_mem_b0_b_119 ), .B (n_3704), .S0 (n_7496), .Y(n_8789));
MX2X1 g34034(.A (u5_mem_b0_b_118 ), .B (n_3707), .S0 (n_7496), .Y(n_8791));
MX2X1 g34037(.A (u5_mem_b0_b_120 ), .B (n_3699), .S0 (n_7496), .Y(n_8787));
MX2X1 g34036(.A (u5_mem_b0_b_92 ), .B (n_3700), .S0 (n_7496), .Y(n_8788));
INVX1 g42580(.A (dma_req_o_b4_b), .Y (n_268));
INVX1 g42581(.A (u11_mem_b0_b_151 ), .Y (n_6357));
INVX1 g41935(.A (n_8182), .Y (n_11036));
INVX1 g42582(.A (u8_wp_b1_b ), .Y (n_178));
NAND2X1 g34244(.A (u8_mem_b3_b_136 ), .B (n_7976), .Y (n_8160));
INVX1 g42587(.A (u9_mem_b0_b_177 ), .Y (n_1724));
OAI21X1 g29907(.A0 (dma_ack_i_b3_b), .A1 (n_118), .B0 (n_11182), .Y(n_11193));
OAI21X1 g29906(.A0 (dma_ack_i_b2_b), .A1 (n_105), .B0 (n_11172), .Y(n_11191));
OAI21X1 g29905(.A0 (dma_ack_i_b1_b), .A1 (n_278), .B0 (n_11183), .Y(n_11194));
OAI21X1 g29904(.A0 (dma_ack_i_b0_b), .A1 (n_271), .B0 (n_11173), .Y(n_11192));
OAI21X1 g29909(.A0 (dma_ack_i_b5_b), .A1 (n_284), .B0 (n_11170), .Y(n_11189));
OAI21X1 g29908(.A0 (dma_ack_i_b4_b), .A1 (n_268), .B0 (n_11171), .Y(n_11190));
NAND2X1 g38815(.A (u4_mem_b3_b_152 ), .B (n_3556), .Y (n_3552));
INVX1 g37108(.A (n_5807), .Y (n_5530));
NAND4X1 g37109(.A (n_11455), .B (n_11456), .C (n_1867), .D (n_2390),.Y (n_5807));
AOI21X1 g38338(.A0 (u5_mem_b3_b_131 ), .A1 (n_5000), .B0 (n_3063), .Y(n_5001));
AOI21X1 g38339(.A0 (u5_mem_b3_b_132 ), .A1 (n_4996), .B0 (n_2929), .Y(n_4999));
INVX1 g37100(.A (n_6769), .Y (n_6070));
NAND4X1 g37101(.A (n_4226), .B (n_2333), .C (n_4123), .D (n_1376), .Y(n_6769));
INVX1 g37102(.A (n_5815), .Y (n_5531));
NAND4X1 g37103(.A (n_11457), .B (n_11458), .C (n_2128), .D (n_1892),.Y (n_5815));
INVX1 g37104(.A (n_11895), .Y (n_5673));
AOI21X1 g38337(.A0 (u5_mem_b3_b ), .A1 (n_5000), .B0 (n_3023), .Y(n_5002));
INVX2 g32887(.A (n_9675), .Y (n_10010));
INVX4 g32885(.A (n_9675), .Y (n_10065));
INVX2 g32882(.A (n_9724), .Y (n_9829));
INVX4 g32883(.A (n_9675), .Y (n_9724));
INVX4 g32880(.A (n_9829), .Y (n_10679));
INVX1 g41932(.A (n_8182), .Y (n_11128));
INVX1 g41875(.A (dma_req_o_b1_b), .Y (n_278));
INVX1 g42830(.A (u9_mem_b1_b_145 ), .Y (n_1727));
INVX1 g42832(.A (u11_mem_b1_b_120 ), .Y (n_6498));
INVX1 g42835(.A (oc4_int_set_715), .Y (n_668));
INVX1 g42836(.A (u10_mem_b1_b_137 ), .Y (n_96));
INVX1 g42837(.A (u10_mem_b1_b_143 ), .Y (n_147));
INVX1 g41933(.A (n_8182), .Y (n_11030));
NOR2X1 g40089(.A (n_2470), .B (n_2691), .Y (n_2142));
NOR2X1 g40088(.A (n_2716), .B (n_1985), .Y (n_2143));
NOR2X1 g40087(.A (n_2144), .B (n_2748), .Y (n_2145));
NOR2X1 g40086(.A (n_821), .B (n_2767), .Y (n_2146));
NOR2X1 g40085(.A (n_945), .B (n_2792), .Y (n_2147));
NOR2X1 g40084(.A (n_2804), .B (n_1985), .Y (n_2149));
NOR2X1 g40083(.A (n_821), .B (n_2720), .Y (n_2151));
NOR2X1 g40081(.A (n_1082), .B (n_2732), .Y (n_2778));
NOR2X1 g40080(.A (n_2786), .B (n_1985), .Y (n_2153));
NOR2X1 g36507(.A (n_829), .B (i4_status), .Y (n_5596));
NAND2X1 g36504(.A (n_1804), .B (n_4081), .Y (n_4082));
NOR2X1 g36503(.A (n_844), .B (i3_status), .Y (n_5597));
NAND2X1 g36502(.A (n_12368), .B (n_6816), .Y (n_6232));
NAND2X1 g36501(.A (n_6816), .B (n_5847), .Y (n_5848));
NAND2X1 g36500(.A (n_12626), .B (n_6816), .Y (n_5850));
AND2X1 g41281(.A (n_710), .B (n_734), .Y (n_841));
INVX1 g41882(.A (u9_mem_b0_b_161 ), .Y (n_6400));
NOR2X1 g36509(.A (n_807), .B (i6_status), .Y (n_5439));
NAND2X1 g36508(.A (n_6781), .B (n_6816), .Y (n_6785));
INVX2 g42956(.A (u5_wp_b0_b ), .Y (n_710));
INVX1 g41883(.A (u9_mem_b3_b_61 ), .Y (n_6912));
AND2X1 g45673(.A (n_782), .B (n_11579), .Y (n_12364));
NAND2X1 g39792(.A (u7_mem_b2_b_43 ), .B (n_12645), .Y (n_2956));
INVX1 g42951(.A (u9_mem_b2_b_88 ), .Y (n_6881));
NAND2X1 g45670(.A (n_12366), .B (u6_mem_b0_b_106 ), .Y (n_12367));
INVX1 g41884(.A (u11_mem_b3_b_71 ), .Y (n_6419));
NAND2X1 g45679(.A (n_12067), .B (n_12375), .Y (n_12376));
INVX1 g41885(.A (u9_mem_b2_b_94 ), .Y (n_6928));
INVX2 g40887(.A (n_1429), .Y (n_3330));
INVX1 g40886(.A (n_3330), .Y (n_2488));
INVX2 g40884(.A (n_1429), .Y (n_3207));
NAND2X2 g40882(.A (n_411), .B (n_705), .Y (n_1226));
INVX2 g40888(.A (n_12614), .Y (n_1429));
INVX1 g36761(.A (o3_status), .Y (n_5398));
INVX1 g36767(.A (o6_status), .Y (n_4070));
INVX1 g36764(.A (o4_status), .Y (n_5396));
INVX1 g42481(.A (n_4088), .Y (n_449));
INVX1 g42482(.A (u9_mem_b0_b_178 ), .Y (n_2500));
INVX1 g42485(.A (u11_mem_b1_b_126 ), .Y (n_6484));
INVX1 g42486(.A (u9_mem_b3_b_59 ), .Y (n_6890));
BUFX3 g41304(.A (n_1059), .Y (n_5480));
INVX4 g40610(.A (wb_din_665), .Y (n_2744));
MX2X1 g38622(.A (u4_mem_b0_b_111 ), .B (wb_din_681), .S0 (n_3765), .Y(n_3777));
NAND2X1 g45557(.A (n_3474), .B (u6_mem_b2_b_38 ), .Y (n_12165));
AOI21X1 g30901(.A0 (n_11631), .A1 (n_11632), .B0 (n_11033), .Y(n_11017));
AOI21X1 g30900(.A0 (n_11639), .A1 (n_11640), .B0 (n_11025), .Y(n_11018));
OAI21X1 g30903(.A0 (n_7295), .A1 (n_7526), .B0 (n_8915), .Y (n_9474));
AOI21X1 g30902(.A0 (n_11641), .A1 (n_11642), .B0 (n_11030), .Y(n_11016));
OAI21X1 g30905(.A0 (n_7387), .A1 (n_8205), .B0 (n_9446), .Y (n_9526));
INVX4 g33303(.A (n_10787), .Y (n_9885));
AND2X1 g30907(.A (n_9691), .B (n_11564), .Y (n_9836));
AND2X1 g30906(.A (n_10338), .B (n_11772), .Y (n_10902));
AND2X1 g30909(.A (n_10337), .B (n_11772), .Y (n_10900));
AND2X1 g30908(.A (n_9961), .B (n_11600), .Y (n_10780));
NAND2X1 g39416(.A (u5_mem_b2_b_31 ), .B (n_12823), .Y (n_11439));
NAND2X1 g39417(.A (n_3259), .B (u5_mem_b0_b_94 ), .Y (n_3192));
NOR2X1 g39410(.A (n_2818), .B (n_1488), .Y (n_1483));
NAND2X1 g39411(.A (u5_mem_b1_b_61 ), .B (n_3236), .Y (n_11444));
NAND2X1 g39412(.A (n_12721), .B (u3_mem_b0_b_107 ), .Y (n_3199));
INVX1 g33309(.A (n_12148), .Y (n_9626));
INVX2 g40617(.A (wb_din_673), .Y (n_2681));
INVX1 g42224(.A (n_9641), .Y (n_685));
INVX1 g42227(.A (u11_mem_b1_b_144 ), .Y (n_1604));
NAND2X1 g34628(.A (u6_mem_b1_b_65 ), .B (n_7758), .Y (n_7797));
OAI21X1 g33909(.A0 (n_4287), .A1 (n_8457), .B0 (n_7613), .Y (n_8936));
NAND2X1 g34624(.A (u6_mem_b1_b_90 ), .B (n_7758), .Y (n_7801));
OAI21X1 g33905(.A0 (n_4412), .A1 (n_8453), .B0 (n_7982), .Y (n_8941));
OAI21X1 g33906(.A0 (n_4329), .A1 (n_8891), .B0 (n_7615), .Y (n_8940));
OAI21X1 g33907(.A0 (n_4288), .A1 (n_8449), .B0 (n_7614), .Y (n_8939));
OAI21X1 g33900(.A0 (n_4885), .A1 (n_8951), .B0 (n_7623), .Y (n_8947));
OAI21X1 g33901(.A0 (n_4956), .A1 (n_8951), .B0 (n_7622), .Y (n_8946));
OAI21X1 g33902(.A0 (n_5146), .A1 (n_8948), .B0 (n_7621), .Y (n_8945));
MX2X1 g31230(.A (n_6027), .B (n_6026), .S0 (n_10839), .Y (n_10834));
MX2X1 g31231(.A (n_6527), .B (n_6526), .S0 (n_10315), .Y (n_10185));
MX2X1 g31232(.A (n_6414), .B (n_6413), .S0 (n_10513), .Y (n_10455));
MX2X1 g31233(.A (n_6416), .B (n_6415), .S0 (n_10137), .Y (n_10184));
MX2X1 g31234(.A (n_6543), .B (n_6542), .S0 (n_10137), .Y (n_10183));
MX2X1 g31235(.A (n_6412), .B (n_6411), .S0 (n_10137), .Y (n_10182));
MX2X1 g31236(.A (n_6525), .B (n_6524), .S0 (n_10513), .Y (n_10454));
MX2X1 g31237(.A (n_6409), .B (n_6408), .S0 (n_10137), .Y (n_10181));
MX2X1 g31238(.A (n_6418), .B (n_6417), .S0 (n_10513), .Y (n_10453));
MX2X1 g31239(.A (n_6407), .B (n_6406), .S0 (n_10315), .Y (n_10180));
INVX1 g42104(.A (n_1198), .Y (n_757));
CLKBUFX1 g42105(.A (n_691), .Y (n_1198));
INVX2 g42106(.A (u8_rp_b1_b ), .Y (n_691));
NAND2X1 g39574(.A (u8_mem_b1_b_65 ), .B (n_12295), .Y (n_11466));
NAND2X1 g39572(.A (n_6042), .B (n_1300), .Y (n_2284));
NAND2X1 g34488(.A (u8_mem_b1_b_60 ), .B (n_7976), .Y (n_7945));
INVX8 g34952(.A (n_7758), .Y (n_7505));
INVX1 g42410(.A (u11_mem_b0_b_154 ), .Y (n_6351));
INVX4 g34485(.A (n_7514), .Y (n_8538));
NAND2X1 g34839(.A (u8_mem_b1_b_61 ), .B (n_7976), .Y (n_7595));
AOI22X1 g35685(.A0 (n_6686), .A1 (i6_dout_644), .B0 (i3_dout_582),.B1 (n_6700), .Y (n_6699));
AOI22X1 g35684(.A0 (n_6686), .A1 (i6_dout_640), .B0 (i3_dout_578),.B1 (n_6700), .Y (n_6702));
AOI22X1 g35687(.A0 (n_6686), .A1 (i6_dout_647), .B0 (i3_dout_585),.B1 (n_6700), .Y (n_6690));
AOI22X1 g35686(.A0 (n_6686), .A1 (i6_dout_646), .B0 (i3_dout_584),.B1 (n_6700), .Y (n_6685));
AOI22X1 g35681(.A0 (n_6686), .A1 (i6_dout), .B0 (i3_dout), .B1(n_6700), .Y (n_6706));
OAI21X1 g35680(.A0 (n_5632), .A1 (u2_res_cnt_b0_b ), .B0 (n_4094), .Y(n_5450));
AOI22X1 g35683(.A0 (n_6686), .A1 (i6_dout_639), .B0 (i3_dout_577),.B1 (n_6700), .Y (n_6703));
AOI22X1 g35682(.A0 (n_6686), .A1 (i6_dout_636), .B0 (i3_dout_574),.B1 (n_6700), .Y (n_6705));
AOI22X1 g35689(.A0 (n_6686), .A1 (i6_dout_651), .B0 (i3_dout_589),.B1 (n_6700), .Y (n_6696));
AOI22X1 g35688(.A0 (n_6686), .A1 (i6_dout_648), .B0 (i3_dout_586),.B1 (n_6700), .Y (n_6697));
NAND2X1 g45527(.A (u4_rp_b0_b ), .B (n_6180), .Y (n_12132));
INVX1 g41967(.A (u11_mem_b0_b_169 ), .Y (n_1634));
INVX1 g41104(.A (n_834), .Y (n_1297));
INVX2 g41966(.A (u4_wp_b0_b ), .Y (n_744));
OAI21X1 g45524(.A0 (n_12135), .A1 (n_12136), .B0 (n_12149), .Y(n_12140));
INVX1 g41965(.A (n_744), .Y (n_1419));
BUFX3 g45879(.A (n_12608), .Y (n_12609));
OAI21X1 g45878(.A0 (n_5571), .A1 (n_6995), .B0 (n_5862), .Y(n_12606));
NAND2X1 g45875(.A (n_6091), .B (n_6241), .Y (n_12602));
NAND2X1 g45874(.A (n_3559), .B (n_5867), .Y (n_12601));
AND2X1 g45877(.A (n_242), .B (n_544), .Y (n_12603));
INVX1 g45876(.A (n_12603), .Y (n_12604));
AOI21X1 g45873(.A0 (n_12601), .A1 (n_12602), .B0 (n_12604), .Y(n_12605));
INVX1 g41962(.A (oc5_int_set_717), .Y (n_611));
INVX1 g40717(.A (n_1176), .Y (n_2135));
INVX1 g41961(.A (u9_mem_b0_b_158 ), .Y (n_6845));
INVX1 g35539(.A (i3_full), .Y (n_632));
INVX4 g40575(.A (wb_din_680), .Y (n_2732));
INVX1 g41960(.A (u11_mem_b0_b_158 ), .Y (n_5947));
NAND4X1 g36888(.A (n_12030), .B (n_3260), .C (n_12031), .D (n_1340),.Y (n_5886));
NAND3X1 g36889(.A (n_576), .B (n_442), .C (n_726), .Y (n_1274));
INVX1 g36882(.A (n_5719), .Y (n_5720));
INVX1 g36880(.A (n_5867), .Y (n_5566));
NAND4X1 g36881(.A (n_11494), .B (n_3270), .C (n_11495), .D (n_1324),.Y (n_5867));
NAND4X1 g36886(.A (n_12034), .B (n_3261), .C (n_12035), .D (n_1544),.Y (n_5857));
INVX1 g36887(.A (n_5886), .Y (n_5564));
NAND4X1 g36884(.A (n_12807), .B (n_12808), .C (n_3268), .D (n_1327),.Y (n_5719));
INVX1 g36885(.A (n_5857), .Y (n_5565));
NAND2X1 g41545(.A (u15_rdd1), .B (u15_crac_rd), .Y (n_414));
OAI21X1 g30723(.A0 (n_5826), .A1 (n_9654), .B0 (n_9653), .Y (n_9655));
OAI21X1 g33430(.A0 (n_5147), .A1 (n_8097), .B0 (n_8069), .Y (n_8436));
INVX1 g41969(.A (oc3_int_set_714), .Y (n_490));
AOI21X1 g38101(.A0 (u8_mem_b2_b_57 ), .A1 (n_4499), .B0 (n_2138), .Y(n_4477));
AOI21X1 g38100(.A0 (u4_mem_b1_b_83 ), .A1 (n_4471), .B0 (n_2115), .Y(n_4478));
AOI21X1 g38103(.A0 (u4_mem_b1_b_75 ), .A1 (n_4507), .B0 (n_2065), .Y(n_4475));
AOI21X1 g38102(.A0 (u6_mem_b2_b_40 ), .A1 (n_4504), .B0 (n_2136), .Y(n_4476));
AOI21X1 g38105(.A0 (u3_mem_b2_b_49 ), .A1 (n_4519), .B0 (n_2191), .Y(n_4474));
AOI21X1 g38104(.A0 (u8_mem_b3_b_147 ), .A1 (n_3879), .B0 (n_1555), .Y(n_3872));
AOI21X1 g38107(.A0 (u8_mem_b3_b_122 ), .A1 (n_3879), .B0 (n_1490), .Y(n_3869));
AOI21X1 g38106(.A0 (u8_mem_b3_b_139 ), .A1 (n_3879), .B0 (n_1272), .Y(n_3871));
AOI21X1 g38109(.A0 (u4_mem_b1_b_70 ), .A1 (n_4471), .B0 (n_2207), .Y(n_4472));
AOI21X1 g38108(.A0 (u4_mem_b1_b ), .A1 (n_4507), .B0 (n_2116), .Y(n_4473));
NOR2X1 g41267(.A (u13_ints_r_b24_b ), .B (ic1_int_set_721), .Y(n_495));
INVX1 g40714(.A (n_1176), .Y (n_2189));
AOI22X1 g37715(.A0 (n_2558), .A1 (n_1244), .B0 (n_5363), .B1(n_1316), .Y (n_1245));
NAND2X1 g39359(.A (u5_mem_b1_b_71 ), .B (n_3236), .Y (n_12796));
INVX1 g42519(.A (dma_req_o_b2_b), .Y (n_105));
NOR2X1 g39358(.A (n_3486), .B (n_2763), .Y (n_3246));
INVX4 g41442(.A (n_982), .Y (n_1488));
NOR2X1 g35308(.A (n_1355), .B (n_12335), .Y (n_7539));
NOR2X1 g40168(.A (n_2686), .B (n_2045), .Y (n_2069));
NOR2X1 g40169(.A (n_2772), .B (n_2067), .Y (n_2068));
NAND2X1 g39356(.A (u5_mem_b2_b_52 ), .B (n_12823), .Y (n_2496));
NOR2X1 g40164(.A (n_2729), .B (n_2008), .Y (n_2073));
NOR2X1 g40165(.A (n_2071), .B (n_2735), .Y (n_2072));
NOR2X1 g40166(.A (n_2085), .B (n_3008), .Y (n_2263));
NOR2X1 g40167(.A (n_2470), .B (n_2684), .Y (n_2070));
NOR2X1 g40160(.A (n_945), .B (n_2741), .Y (n_2079));
NOR2X1 g40161(.A (n_935), .B (n_2744), .Y (n_2077));
NOR2X1 g40162(.A (n_2120), .B (n_2716), .Y (n_2075));
NOR2X1 g40163(.A (n_2470), .B (n_2763), .Y (n_2074));
INVX1 g42518(.A (oc5_cfg_1019), .Y (n_469));
INVX1 g40712(.A (n_1176), .Y (n_2218));
NAND2X1 g39879(.A (n_12679), .B (u5_mem_b0_b_113 ), .Y (n_3846));
NAND2X1 g45558(.A (n_2419), .B (u6_mem_b3_b_131 ), .Y (n_12166));
NAND4X1 g37593(.A (u26_ps_cnt_b3_b ), .B (u26_ps_cnt_b1_b ), .C(u26_ps_cnt_b0_b ), .D (n_681), .Y (n_1775));
AND2X1 g37592(.A (n_3549), .B (n_4633), .Y (n_4634));
AOI21X1 g37591(.A0 (n_5225), .A1 (n_675), .B0 (wb_addr_i_b6_b), .Y(n_2608));
NAND3X1 g37590(.A (n_581), .B (n_1006), .C (u12_re1), .Y (n_1815));
NOR2X1 g37597(.A (n_1209), .B (n_2368), .Y (n_2570));
NOR2X1 g37596(.A (n_1199), .B (n_2302), .Y (n_3941));
AND2X1 g37595(.A (n_2371), .B (n_3942), .Y (n_3943));
AOI21X1 g38412(.A0 (u6_mem_b1_b_74 ), .A1 (n_5112), .B0 (n_2683), .Y(n_4941));
NOR2X1 g37599(.A (n_1224), .B (n_2513), .Y (n_2569));
AOI21X1 g38147(.A0 (u4_mem_b2_b_42 ), .A1 (n_4439), .B0 (n_2111), .Y(n_4436));
OAI21X1 g33683(.A0 (n_4983), .A1 (n_9290), .B0 (n_7856), .Y (n_9218));
OAI21X1 g33682(.A0 (n_4984), .A1 (n_9290), .B0 (n_7857), .Y (n_9219));
OAI21X1 g33681(.A0 (n_4985), .A1 (n_9290), .B0 (n_7858), .Y (n_9221));
OAI21X1 g33680(.A0 (n_4986), .A1 (n_9290), .B0 (n_7859), .Y (n_9222));
OAI21X1 g33687(.A0 (n_4979), .A1 (n_9212), .B0 (n_7852), .Y (n_9213));
OAI21X1 g33686(.A0 (n_4980), .A1 (n_9212), .B0 (n_7853), .Y (n_9214));
OAI21X1 g33685(.A0 (n_4981), .A1 (n_9230), .B0 (n_7854), .Y (n_9216));
OAI21X1 g33684(.A0 (n_4982), .A1 (n_9230), .B0 (n_7855), .Y (n_9217));
AOI21X1 g38141(.A0 (u4_mem_b1_b_67 ), .A1 (n_4471), .B0 (n_1958), .Y(n_4444));
OAI21X1 g33689(.A0 (n_4977), .A1 (n_9212), .B0 (n_7850), .Y (n_9210));
NAND2X1 g38972(.A (u8_mem_b3_b_148 ), .B (n_2468), .Y (n_2389));
AOI21X1 g38140(.A0 (u4_mem_b1_b_66 ), .A1 (n_4471), .B0 (n_1940), .Y(n_4445));
AOI21X1 g38414(.A0 (u6_mem_b1_b_83 ), .A1 (n_5112), .B0 (n_2817), .Y(n_4940));
AOI22X1 g37661(.A0 (in_slt_413), .A1 (n_1406), .B0 (in_slt_415), .B1(n_4624), .Y (n_4625));
AOI22X1 g37663(.A0 (in_slt_397), .A1 (n_1406), .B0 (u9_din_tmp_42),.B1 (n_2368), .Y (n_4621));
OAI21X1 g37379(.A0 (u9_mem_b0_b_180 ), .A1 (n_6856), .B0 (n_4647), .Y(n_5487));
OAI21X1 g37378(.A0 (u10_mem_b0_b_169 ), .A1 (n_6341), .B0 (n_5240), .Y(n_5665));
OAI21X1 g37377(.A0 (u11_mem_b0_b_173 ), .A1 (n_6359), .B0 (n_5239), .Y(n_5666));
AOI22X1 g37376(.A0 (n_5272), .A1 (u13_intm_r_b14_b ), .B0 (n_5277),.B1 (crac_din_705), .Y (n_5251));
AOI22X1 g37375(.A0 (n_5277), .A1 (crac_out_862), .B0 (n_6972), .B1(oc2_cfg_984), .Y (n_3983));
INVX1 g37374(.A (n_3983), .Y (n_4681));
AOI22X1 g37373(.A0 (n_5591), .A1 (n_4683), .B0 (n_6972), .B1(oc2_cfg_985), .Y (n_4685));
NAND2X1 g38812(.A (u4_mem_b3_b_138 ), .B (n_4258), .Y (n_4261));
AOI22X1 g37370(.A0 (n_5272), .A1 (u13_intm_r_b19_b ), .B0(u13_ints_r_b19_b ), .B1 (n_4726), .Y (n_4686));
NAND2X1 g39752(.A (n_12389), .B (u4_mem_b0_b_97 ), .Y (n_11658));
AOI22X1 g37666(.A0 (in_slt_398), .A1 (n_1406), .B0 (u9_din_tmp_43),.B1 (n_2368), .Y (n_4619));
INVX8 g41566(.A (n_1448), .Y (n_3089));
INVX2 g41175(.A (n_1299), .Y (n_3415));
NOR2X1 g39756(.A (n_4996), .B (n_2707), .Y (n_2975));
NOR2X1 g39754(.A (n_4961), .B (n_2831), .Y (n_2976));
INVX8 g41040(.A (n_1027), .Y (n_2470));
NAND2X1 g39758(.A (n_2325), .B (in_slt_446), .Y (n_2252));
NAND2X1 g41042(.A (u4_wp_b0_b ), .B (n_444), .Y (n_821));
NAND2X1 g38976(.A (u7_mem_b3_b_132 ), .B (n_1538), .Y (n_1383));
INVX1 g41043(.A (n_1412), .Y (n_3257));
INVX1 g41177(.A (n_1049), .Y (n_1299));
NAND2X1 g32627(.A (u9_wp_b2_b ), .B (n_9514), .Y (n_9687));
NAND2X1 g38977(.A (u8_mem_b3_b_152 ), .B (n_2468), .Y (n_2385));
CLKBUFX1 g41178(.A (n_1049), .Y (n_4624));
MX2X1 g38626(.A (u4_mem_b0_b_115 ), .B (wb_din_685), .S0 (n_835), .Y(n_3768));
INVX1 g42510(.A (n_551), .Y (n_761));
INVX8 g35056(.A (o4_we), .Y (n_7984));
NAND2X1 g38978(.A (u7_mem_b3_b_150 ), .B (n_1546), .Y (n_1386));
INVX2 g42039(.A (n_5772), .Y (n_6318));
INVX1 g42030(.A (u10_mem_b0_b_180 ), .Y (n_1864));
NOR2X1 g40196(.A (n_2775), .B (n_2763), .Y (n_2723));
OAI21X1 g35946(.A0 (n_5684), .A1 (n_7077), .B0 (n_6158), .Y (n_7055));
OAI21X1 g35947(.A0 (n_5669), .A1 (n_7063), .B0 (n_5801), .Y (n_7054));
OAI21X1 g35944(.A0 (n_5546), .A1 (n_6981), .B0 (n_5806), .Y (n_6978));
OAI21X1 g35945(.A0 (n_5700), .A1 (n_7077), .B0 (n_6162), .Y (n_7056));
OAI21X1 g35942(.A0 (n_5673), .A1 (n_7077), .B0 (n_6164), .Y (n_7058));
OAI21X1 g35943(.A0 (n_5672), .A1 (n_7063), .B0 (n_6221), .Y (n_7057));
OAI21X1 g35940(.A0 (n_5537), .A1 (n_7063), .B0 (n_5824), .Y (n_6979));
INVX1 g35233(.A (n_7396), .Y (n_8894));
NAND2X1 g40769(.A (n_746), .B (u7_wp_b1_b ), .Y (n_938));
INVX1 g35238(.A (n_7396), .Y (n_8891));
INVX1 g35239(.A (n_7396), .Y (n_8933));
OAI21X1 g35948(.A0 (n_5721), .A1 (n_7063), .B0 (n_5894), .Y (n_7053));
INVX1 g40718(.A (n_1176), .Y (n_2081));
INVX1 g41913(.A (u11_mem_b3_b_61 ), .Y (n_6556));
OR2X1 g39198(.A (n_7120), .B (n_2567), .Y (n_2300));
NAND2X1 g39195(.A (n_12840), .B (u4_mem_b0_b_93 ), .Y (n_3388));
NAND2X1 g39194(.A (n_3252), .B (u7_mem_b0_b_116 ), .Y (n_3389));
NAND2X1 g39196(.A (u4_mem_b2_b_31 ), .B (n_12079), .Y (n_2304));
NOR2X1 g39191(.A (n_5138), .B (n_2794), .Y (n_3391));
NOR2X1 g39190(.A (n_3089), .B (n_2864), .Y (n_3392));
NAND3X1 g39193(.A (u4_mem_b0_b_92 ), .B (n_868), .C (n_1923), .Y(n_1491));
NAND2X1 g39192(.A (n_11798), .B (u8_mem_b0_b_102 ), .Y (n_11453));
NAND2X1 g38837(.A (u7_mem_b3_b_146 ), .B (n_1546), .Y (n_1547));
MX2X1 g38627(.A (u4_mem_b0_b_116 ), .B (wb_din_686), .S0 (n_3765), .Y(n_3766));
NAND2X1 g38836(.A (u5_mem_b3_b_133 ), .B (n_1543), .Y (n_1325));
MX2X1 g34013(.A (u3_mem_b0_b_116 ), .B (n_3586), .S0 (n_8700), .Y(n_8810));
MX2X1 g34012(.A (u4_mem_b0_b_99 ), .B (n_3752), .S0 (n_7499), .Y(n_9430));
NAND2X1 g34547(.A (u5_mem_b2_b_59 ), .B (n_7870), .Y (n_7880));
NAND2X1 g34546(.A (u5_mem_b2_b_58 ), .B (n_7870), .Y (n_7881));
MX2X1 g34017(.A (u5_mem_b0_b_102 ), .B (n_3735), .S0 (n_7496), .Y(n_8806));
MX2X1 g34016(.A (u5_mem_b0_b_101 ), .B (n_3737), .S0 (n_7496), .Y(n_8807));
MX2X1 g34015(.A (u5_mem_b0_b_100 ), .B (n_3739), .S0 (n_7496), .Y(n_8808));
MX2X1 g34019(.A (u5_mem_b0_b_104 ), .B (n_3734), .S0 (n_7496), .Y(n_9428));
MX2X1 g34018(.A (u5_mem_b0_b_103 ), .B (n_3624), .S0 (n_7496), .Y(n_9429));
NAND2X1 g34549(.A (u5_mem_b2_b_32 ), .B (n_7870), .Y (n_7878));
NAND2X1 g34548(.A (u5_mem_b2_b_31 ), .B (n_7870), .Y (n_7879));
NAND2X1 g38831(.A (u6_mem_b3_b_132 ), .B (n_2419), .Y (n_2447));
INVX1 g43071(.A (u10_mem_b1_b_123 ), .Y (n_6411));
INVX1 g43070(.A (u11_mem_b0_b_177 ), .Y (n_1596));
AOI21X1 g37691(.A0 (n_6585), .A1 (n_1316), .B0 (n_2346), .Y (n_3929));
NAND2X1 g39771(.A (u8_mem_b2_b_53 ), .B (n_2366), .Y (n_2301));
NAND2X1 g38833(.A (n_9641), .B (n_1889), .Y (n_3549));
NAND2X1 g45559(.A (n_12169), .B (u6_mem_b1_b_69 ), .Y (n_12170));
NAND2X2 g40869(.A (n_744), .B (u4_wp_b1_b ), .Y (n_935));
NOR2X1 g45539(.A (oc1_cfg_975), .B (oc1_cfg_976), .Y (n_12144));
INVX1 g40868(.A (n_935), .Y (n_1019));
INVX1 g40713(.A (n_1176), .Y (n_2154));
OAI21X1 g33578(.A0 (n_5096), .A1 (n_9349), .B0 (n_7975), .Y (n_9350));
INVX2 g45624(.A (n_12303), .Y (n_12301));
INVX1 g42852(.A (u10_mem_b2_b_116 ), .Y (n_42));
INVX1 g42850(.A (n_434), .Y (n_4738));
INVX1 g42851(.A (ic1_cfg_1035), .Y (n_434));
INVX1 g42856(.A (u9_mem_b1_b_127 ), .Y (n_6937));
NAND2X1 g37163(.A (n_3908), .B (n_2273), .Y (n_6521));
NAND2X1 g37160(.A (n_4614), .B (n_3515), .Y (n_6927));
NAND2X1 g37161(.A (n_3909), .B (n_1795), .Y (n_6592));
NAND2X1 g37166(.A (n_3903), .B (n_1564), .Y (n_6514));
NAND2X1 g37167(.A (n_3902), .B (n_2227), .Y (n_6510));
NAND2X1 g37164(.A (n_3907), .B (n_2269), .Y (n_6478));
NAND2X1 g37165(.A (n_3904), .B (n_2345), .Y (n_6586));
NAND2X1 g37168(.A (n_2520), .B (n_2268), .Y (n_6014));
NAND2X1 g37169(.A (n_3900), .B (n_2288), .Y (n_6465));
AOI21X1 g38318(.A0 (u5_mem_b2_b_50 ), .A1 (n_4370), .B0 (n_2040), .Y(n_4364));
AOI21X1 g38319(.A0 (u6_mem_b1_b_82 ), .A1 (n_5112), .B0 (n_2650), .Y(n_5007));
NAND2X1 g36564(.A (n_5818), .B (n_6201), .Y (n_5817));
NAND2X1 g36567(.A (n_6765), .B (n_784), .Y (n_6766));
NAND2X1 g36566(.A (n_11855), .B (n_6201), .Y (n_6197));
NAND2X1 g36569(.A (n_6194), .B (n_12115), .Y (n_6195));
NAND2X1 g36568(.A (n_2615), .B (u2_to_cnt_b5_b ), .Y (n_2616));
INVX1 g42931(.A (u11_mem_b2_b_100 ), .Y (n_461));
INVX1 g42932(.A (u10_mem_b2_b_109 ), .Y (n_2556));
INVX2 g45614(.A (u8_rp_b2_b ), .Y (n_12281));
INVX1 g42937(.A (oc1_cfg_979), .Y (n_510));
INVX1 g42939(.A (u10_mem_b1_b_134 ), .Y (n_5974));
INVX1 g42938(.A (u9_mem_b0_b_173 ), .Y (n_1733));
INVX1 g45626(.A (n_637), .Y (n_12304));
NAND2X1 g37710(.A (n_2425), .B (n_3080), .Y (n_12051));
NAND2X1 g36789(.A (n_1639), .B (n_1698), .Y (n_4062));
NAND2X1 g36788(.A (n_1860), .B (n_1761), .Y (n_4063));
NAND2X1 g36785(.A (n_1697), .B (n_1848), .Y (n_4066));
NAND2X1 g36784(.A (n_1770), .B (n_1768), .Y (n_4067));
NAND2X1 g36786(.A (n_1765), .B (n_1764), .Y (n_4065));
INVX1 g36781(.A (n_6765), .Y (n_6085));
AND2X1 g36780(.A (n_1553), .B (n_1819), .Y (n_1276));
NAND2X1 g36783(.A (n_825), .B (n_2513), .Y (n_1816));
NAND4X1 g36782(.A (n_3509), .B (n_3056), .C (n_4249), .D (n_2420), .Y(n_6765));
INVX1 g42049(.A (u10_mem_b0_b_178 ), .Y (n_2539));
INVX4 g45620(.A (n_12303), .Y (n_12291));
AOI22X1 g37786(.A0 (n_5994), .A1 (n_1575), .B0 (n_6023), .B1(n_1831), .Y (n_1655));
AOI22X1 g37787(.A0 (n_6542), .A1 (n_2530), .B0 (n_6630), .B1(n_2534), .Y (n_2531));
AOI22X1 g37784(.A0 (n_2558), .A1 (n_6339), .B0 (n_6575), .B1(n_1316), .Y (n_1237));
AOI22X1 g37785(.A0 (n_1756), .A1 (n_5953), .B0 (n_5990), .B1(n_1643), .Y (n_1656));
NAND2X1 g37782(.A (n_2403), .B (n_3038), .Y (n_12061));
AOI22X1 g37783(.A0 (in_slt_401), .A1 (n_1406), .B0 (u9_din_tmp_46),.B1 (n_2368), .Y (n_4584));
AOI22X1 g37780(.A0 (n_6460), .A1 (n_1575), .B0 (n_6419), .B1(n_1831), .Y (n_1658));
AOI22X1 g37781(.A0 (n_2558), .A1 (n_6382), .B0 (n_6463), .B1(n_1839), .Y (n_1657));
AOI22X1 g37788(.A0 (n_1756), .A1 (n_5951), .B0 (n_5988), .B1(n_1643), .Y (n_1654));
AOI22X1 g37789(.A0 (n_6479), .A1 (n_1575), .B0 (n_6428), .B1(n_1831), .Y (n_1653));
MX2X1 g33096(.A (n_227), .B (wb_din_661), .S0 (n_8643), .Y (n_8646));
MX2X1 g33097(.A (n_306), .B (wb_din_662), .S0 (n_8643), .Y (n_8644));
MX2X1 g33094(.A (n_177), .B (wb_din_674), .S0 (n_8643), .Y (n_8649));
MX2X1 g33095(.A (n_170), .B (wb_din_675), .S0 (n_8643), .Y (n_8648));
MX2X1 g33092(.A (n_338), .B (wb_din_672), .S0 (n_8643), .Y (n_8652));
MX2X1 g33093(.A (n_179), .B (wb_din_673), .S0 (n_8643), .Y (n_8651));
MX2X1 g33091(.A (n_138), .B (wb_din_671), .S0 (n_8643), .Y (n_8653));
MX2X1 g33098(.A (n_130), .B (wb_din_664), .S0 (n_8643), .Y (n_8642));
OAI21X1 g31780(.A0 (n_4848), .A1 (n_9631), .B0 (n_9835), .Y(n_10340));
AOI21X1 g31781(.A0 (n_1549), .A1 (n_12303), .B0 (n_11894), .Y(n_9966));
AOI21X1 g31782(.A0 (n_2488), .A1 (n_1918), .B0 (n_12339), .Y(n_9965));
OAI21X1 g31783(.A0 (n_4850), .A1 (n_9514), .B0 (n_9687), .Y (n_9841));
AOI21X1 g31784(.A0 (n_10790), .A1 (n_10787), .B0 (n_9941), .Y(n_10791));
AOI21X1 g31785(.A0 (n_10788), .A1 (n_10787), .B0 (n_9940), .Y(n_10789));
OAI21X1 g31038(.A0 (n_5337), .A1 (n_10820), .B0 (n_10371), .Y(n_10875));
AOI21X1 g31787(.A0 (n_10785), .A1 (n_9931), .B0 (n_9921), .Y(n_10786));
AOI21X1 g31788(.A0 (n_10783), .A1 (n_9931), .B0 (n_9920), .Y(n_10784));
OAI21X1 g31037(.A0 (n_5411), .A1 (n_10880), .B0 (n_10372), .Y(n_10876));
OAI21X1 g31034(.A0 (n_5338), .A1 (n_10880), .B0 (n_10375), .Y(n_10881));
OAI21X1 g31035(.A0 (n_5381), .A1 (n_10880), .B0 (n_10374), .Y(n_10879));
OAI21X1 g31032(.A0 (n_5320), .A1 (n_10820), .B0 (n_10378), .Y(n_10884));
OAI21X1 g31033(.A0 (n_5325), .A1 (n_10820), .B0 (n_10377), .Y(n_10882));
OAI21X1 g31030(.A0 (n_5326), .A1 (n_10880), .B0 (n_10380), .Y(n_10886));
OAI21X1 g31031(.A0 (n_5319), .A1 (n_10820), .B0 (n_10379), .Y(n_10885));
OAI21X1 g33469(.A0 (n_4511), .A1 (n_8440), .B0 (n_8105), .Y (n_8390));
OAI21X1 g33468(.A0 (n_4517), .A1 (n_8393), .B0 (n_8106), .Y (n_8391));
INVX1 g33320(.A (n_12607), .Y (n_11491));
NAND2X1 g34307(.A (u3_mem_b3_b_141 ), .B (n_8101), .Y (n_8089));
NOR2X1 g30929(.A (n_9487), .B (n_9589), .Y (n_9590));
NOR2X1 g30928(.A (n_9549), .B (n_9647), .Y (n_9648));
INVX4 g33324(.A (n_10518), .Y (n_10645));
INVX2 g41006(.A (n_1416), .Y (n_2775));
INVX8 g33327(.A (n_9876), .Y (n_10518));
NOR2X1 g30923(.A (n_4827), .B (n_9597), .Y (n_9593));
NOR2X1 g30922(.A (n_3994), .B (n_9597), .Y (n_9594));
NOR2X1 g30921(.A (n_2630), .B (n_9597), .Y (n_9595));
NOR2X1 g30920(.A (n_3849), .B (n_9597), .Y (n_9596));
NOR2X1 g30927(.A (n_9489), .B (n_9591), .Y (n_9592));
NAND2X1 g30926(.A (n_9844), .B (n_9831), .Y (n_10333));
NAND2X1 g30925(.A (n_9759), .B (n_9734), .Y (n_9951));
NAND2X1 g30924(.A (n_10086), .B (n_9910), .Y (n_10777));
NAND2X1 g34304(.A (u3_mem_b3_b_140 ), .B (n_8101), .Y (n_8091));
AOI22X1 g37713(.A0 (u9_din_tmp_52), .A1 (n_2368), .B0 (in_slt_409),.B1 (n_4624), .Y (n_2561));
INVX1 g42207(.A (oc2_cfg_985), .Y (n_544));
NAND2X1 g34303(.A (u3_mem_b3_b_139 ), .B (n_8101), .Y (n_8092));
INVX1 g42205(.A (u10_mem_b1_b_138 ), .Y (n_90));
INVX1 g42204(.A (oc0_int_set_708), .Y (n_492));
INVX1 g42202(.A (n_5788), .Y (n_802));
NAND2X1 g34302(.A (u3_mem_b3_b_138 ), .B (n_8097), .Y (n_8093));
MX2X1 g31258(.A (n_5484), .B (n_1680), .S0 (n_10303), .Y (n_10163));
MX2X1 g31259(.A (n_5468), .B (n_1738), .S0 (n_10303), .Y (n_10162));
OAI21X1 g33461(.A0 (n_4392), .A1 (n_8393), .B0 (n_8115), .Y (n_8399));
MX2X1 g31252(.A (n_6399), .B (n_6398), .S0 (n_10235), .Y (n_10169));
MX2X1 g31253(.A (n_6397), .B (n_6396), .S0 (n_10235), .Y (n_10168));
MX2X1 g31250(.A (n_6401), .B (n_6400), .S0 (n_10250), .Y (n_10172));
MX2X1 g31251(.A (n_6393), .B (n_6392), .S0 (n_10250), .Y (n_10170));
MX2X1 g31256(.A (n_6863), .B (n_6862), .S0 (n_10250), .Y (n_10165));
MX2X1 g31257(.A (n_5486), .B (n_1742), .S0 (n_10250), .Y (n_10164));
MX2X1 g31254(.A (n_6867), .B (n_6866), .S0 (n_10303), .Y (n_10167));
MX2X1 g31255(.A (n_6865), .B (n_6864), .S0 (n_10303), .Y (n_10166));
NOR2X1 g39692(.A (n_2772), .B (n_1488), .Y (n_1477));
NOR2X1 g39693(.A (n_3117), .B (n_2864), .Y (n_3018));
NAND2X1 g39690(.A (u3_mem_b2_b_43 ), .B (n_3207), .Y (n_3019));
NOR2X1 g39696(.A (n_3453), .B (n_2864), .Y (n_3015));
NAND2X1 g39697(.A (u3_mem_b1_b_65 ), .B (n_3316), .Y (n_3014));
NAND2X1 g39694(.A (u8_mem_b1_b_89 ), .B (n_12291), .Y (n_3016));
NAND2X1 g39695(.A (u7_mem_b2_b_55 ), .B (n_12650), .Y (n_4142));
NAND2X1 g39699(.A (n_11789), .B (u8_mem_b0_b_94 ), .Y (n_11463));
INVX1 g41893(.A (u10_mem_b0_b_151 ), .Y (n_6342));
INVX2 g45857(.A (u5_rp_b2_b ), .Y (n_12581));
AOI22X1 g37644(.A0 (n_2502), .A1 (n_6859), .B0 (n_6879), .B1(n_1859), .Y (n_1719));
INVX1 g39036(.A (n_4778), .Y (n_3492));
NAND2X1 g39034(.A (u4_mem_b1_b_67 ), .B (n_12272), .Y (n_11661));
NAND2X1 g39035(.A (u4_mem_b2_b_57 ), .B (n_12091), .Y (n_3493));
NAND2X1 g39032(.A (u3_mem_b2_b_57 ), .B (n_3330), .Y (n_3495));
NAND2X1 g39033(.A (u6_mem_b2_b_57 ), .B (n_3423), .Y (n_3494));
NAND2X1 g39030(.A (u4_mem_b2_b_54 ), .B (n_12079), .Y (n_3497));
NAND2X1 g39031(.A (u4_mem_b1_b_76 ), .B (n_12259), .Y (n_4243));
AOI22X1 g37712(.A0 (n_2558), .A1 (n_1246), .B0 (n_5520), .B1(n_1316), .Y (n_1247));
NAND3X1 g39038(.A (u6_mem_b0_b_91 ), .B (n_888), .C (n_11585), .Y(n_1415));
NAND2X1 g39039(.A (u7_mem_b1_b_82 ), .B (n_4130), .Y (n_4240));
INVX1 g42534(.A (u9_mem_b1_b_130 ), .Y (n_6540));
AOI21X1 g30071(.A0 (n_10397), .A1 (n_11002), .B0 (n_5839), .Y(n_11162));
AOI21X1 g30070(.A0 (n_11512), .A1 (n_11513), .B0 (n_12585), .Y(n_11163));
AND2X1 g30073(.A (n_10968), .B (n_9833), .Y (n_11152));
AND2X1 g30072(.A (n_10969), .B (n_991), .Y (n_11153));
AOI21X1 g30075(.A0 (n_11508), .A1 (n_11509), .B0 (n_11144), .Y(n_11160));
AOI21X1 g30074(.A0 (n_11510), .A1 (n_11511), .B0 (n_1870), .Y(n_11161));
OAI21X1 g30077(.A0 (n_5942), .A1 (n_10985), .B0 (n_10986), .Y(n_11150));
OAI21X1 g30076(.A0 (n_6328), .A1 (n_10992), .B0 (n_10993), .Y(n_11151));
INVX1 g42535(.A (u9_mem_b3_b_79 ), .Y (n_5372));
INVX4 g34977(.A (n_8141), .Y (n_8700));
INVX1 g45581(.A (n_12823), .Y (n_12214));
INVX2 g32780(.A (n_9633), .Y (n_10024));
INVX4 g32783(.A (n_9737), .Y (n_10308));
NAND2X1 g39254(.A (n_12204), .B (u6_mem_b0_b_103 ), .Y (n_11699));
INVX4 g32787(.A (n_9737), .Y (n_10045));
INVX2 g41524(.A (n_638), .Y (n_1316));
AOI21X1 g38129(.A0 (u3_mem_b1_b_84 ), .A1 (n_5157), .B0 (n_2833), .Y(n_5116));
AOI21X1 g38128(.A0 (u4_mem_b1_b_85 ), .A1 (n_4507), .B0 (n_1962), .Y(n_4454));
AOI21X1 g38123(.A0 (u7_mem_b1_b_63 ), .A1 (n_5118), .B0 (n_2738), .Y(n_5117));
AOI21X1 g38122(.A0 (u4_mem_b1_b_80 ), .A1 (n_4507), .B0 (n_2063), .Y(n_4459));
AOI21X1 g38121(.A0 (u4_mem_b1_b_79 ), .A1 (n_4471), .B0 (n_2208), .Y(n_4460));
AOI21X1 g38120(.A0 (u4_mem_b1_b_60 ), .A1 (n_4507), .B0 (n_2184), .Y(n_4461));
AOI21X1 g38127(.A0 (u4_mem_b1_b_84 ), .A1 (n_4471), .B0 (n_2113), .Y(n_4455));
AOI21X1 g38126(.A0 (u4_mem_b1_b_82 ), .A1 (n_4471), .B0 (n_2070), .Y(n_4456));
AOI21X1 g38125(.A0 (u6_mem_b2_b_32 ), .A1 (n_4544), .B0 (n_2094), .Y(n_4457));
AOI21X1 g38124(.A0 (u4_mem_b1_b_81 ), .A1 (n_4471), .B0 (n_2061), .Y(n_4458));
INVX1 g42614(.A (u9_mem_b1_b_143 ), .Y (n_45));
NAND2X1 g45933(.A (n_3209), .B (u5_mem_b1_b_77 ), .Y (n_12674));
NAND2X1 g45935(.A (n_1543), .B (u5_mem_b3_b_139 ), .Y (n_12676));
INVX1 g41862(.A (u9_mem_b3_b_65 ), .Y (n_6905));
INVX1 g42536(.A (u9_mem_b0_b_172 ), .Y (n_1562));
AOI22X1 g37804(.A0 (n_6408), .A1 (n_2530), .B0 (n_6612), .B1(n_2544), .Y (n_2529));
CLKBUFX3 g41529(.A (n_1084), .Y (n_2330));
NAND2X1 g45939(.A (n_12583), .B (n_12581), .Y (n_12677));
NAND2X1 g41528(.A (u10_rp_b1_b ), .B (u10_rp_b0_b ), .Y (n_638));
INVX1 g41867(.A (u10_mem_b1_b_141 ), .Y (n_232));
OAI21X1 g33526(.A0 (n_4453), .A1 (n_9333), .B0 (n_8031), .Y (n_8320));
OAI21X1 g33527(.A0 (n_4508), .A1 (n_8318), .B0 (n_8030), .Y (n_8319));
OAI21X1 g33524(.A0 (n_4455), .A1 (n_8318), .B0 (n_8033), .Y (n_8322));
OAI21X1 g33525(.A0 (n_4454), .A1 (n_8333), .B0 (n_8032), .Y (n_8321));
OAI21X1 g33522(.A0 (n_4456), .A1 (n_9349), .B0 (n_8035), .Y (n_8325));
OAI21X1 g33523(.A0 (n_4478), .A1 (n_9349), .B0 (n_8034), .Y (n_8324));
OAI21X1 g33520(.A0 (n_4459), .A1 (n_8333), .B0 (n_8037), .Y (n_8327));
OAI21X1 g33521(.A0 (n_4458), .A1 (n_9349), .B0 (n_8036), .Y (n_8326));
OAI21X1 g33528(.A0 (n_4514), .A1 (n_9333), .B0 (n_8029), .Y (n_8317));
NAND2X1 g45813(.A (u4_mem_b1_b_63 ), .B (n_12252), .Y (n_12527));
NAND4X1 g45811(.A (n_12526), .B (n_12527), .C (n_12528), .D(n_12529), .Y (n_12530));
INVX1 g41869(.A (u9_mem_b2_b_113 ), .Y (n_365));
NOR2X1 g45816(.A (oc1_cfg_975), .B (n_283), .Y (n_12531));
NAND2X1 g38789(.A (u8_mem_b3_b_151 ), .B (n_2468), .Y (n_2469));
INVX2 g37575(.A (n_5629), .Y (n_5630));
AOI22X1 g38786(.A0 (n_4253), .A1 (n_784), .B0 (n_6821), .B1 (n_762),.Y (n_4854));
AOI22X1 g38785(.A0 (n_3522), .A1 (u7_rp_b0_b ), .B0 (n_12634), .B1(n_754), .Y (n_4266));
OAI21X1 g38784(.A0 (n_1412), .A1 (n_3559), .B0 (n_923), .Y (n_3560));
NAND2X1 g37571(.A (n_5645), .B (n_4153), .Y (n_5229));
NOR2X1 g37570(.A (n_5307), .B (n_6649), .Y (n_4640));
INVX1 g38780(.A (n_4104), .Y (n_3561));
OAI21X1 g33669(.A0 (n_5001), .A1 (n_9235), .B0 (n_7871), .Y (n_9236));
OAI21X1 g33668(.A0 (n_5002), .A1 (n_9235), .B0 (n_7872), .Y (n_9237));
OAI21X1 g33665(.A0 (n_4353), .A1 (n_9264), .B0 (n_7875), .Y (n_9240));
OAI21X1 g33664(.A0 (n_4354), .A1 (n_9202), .B0 (n_7876), .Y (n_9241));
OAI21X1 g33667(.A0 (n_4351), .A1 (n_9307), .B0 (n_7873), .Y (n_9238));
OAI21X1 g33666(.A0 (n_4352), .A1 (n_9264), .B0 (n_7874), .Y (n_9239));
OAI21X1 g33661(.A0 (n_4355), .A1 (n_9286), .B0 (n_7879), .Y (n_9244));
OAI21X1 g33660(.A0 (n_4356), .A1 (n_9235), .B0 (n_7880), .Y (n_9245));
OAI21X1 g33663(.A0 (n_4308), .A1 (n_9202), .B0 (n_7877), .Y (n_9242));
OAI21X1 g33662(.A0 (n_4306), .A1 (n_9212), .B0 (n_7878), .Y (n_9243));
NOR2X1 g39079(.A (n_5138), .B (n_2831), .Y (n_3467));
MX2X1 g31809(.A (n_4074), .B (n_4075), .S0 (n_9690), .Y (n_9691));
MX2X1 g31808(.A (u11_wp_b1_b ), .B (n_4073), .S0 (n_9672), .Y(n_10338));
AOI22X1 g31807(.A0 (n_9795), .A1 (u15_crac_rd), .B0 (crac_out_876),.B1 (u15_crac_we_r), .Y (n_10781));
INVX1 g31806(.A (n_10781), .Y (n_10903));
AOI21X1 g31805(.A0 (n_9952), .A1 (n_9873), .B0 (n_10573), .Y(n_10973));
AOI21X1 g31804(.A0 (n_9602), .A1 (n_9873), .B0 (n_10574), .Y(n_10974));
AOI21X1 g31803(.A0 (n_10976), .A1 (n_10605), .B0 (n_10587), .Y(n_10977));
AOI21X1 g31802(.A0 (n_10978), .A1 (n_10605), .B0 (n_10589), .Y(n_10979));
AOI21X1 g31801(.A0 (n_12656), .A1 (n_1907), .B0 (n_11890), .Y(n_9962));
AOI21X1 g31800(.A0 (n_10981), .A1 (n_10617), .B0 (n_10613), .Y(n_10982));
NOR2X1 g39957(.A (n_2735), .B (n_1488), .Y (n_1457));
NOR2X1 g40376(.A (n_2705), .B (n_2684), .Y (n_2649));
AOI22X1 g37319(.A0 (n_4729), .A1 (n_8197), .B0 (n_5591), .B1(n_4734), .Y (n_4735));
AOI21X1 g31400(.A0 (n_11889), .A1 (n_1184), .B0 (n_9989), .Y(n_10402));
INVX1 g39073(.A (n_4757), .Y (n_3470));
MX2X1 g37310(.A (u10_mem_b1_b_142 ), .B (n_5287), .S0 (n_6475), .Y(n_5288));
MX2X1 g37313(.A (u9_mem_b2_b_114 ), .B (n_4743), .S0 (n_5732), .Y(n_4744));
MX2X1 g37312(.A (u10_mem_b2_b_110 ), .B (n_5282), .S0 (n_5424), .Y(n_5283));
AOI22X1 g37315(.A0 (n_4729), .A1 (n_1481), .B0 (n_5591), .B1(n_11564), .Y (n_4742));
MX2X1 g37314(.A (u11_mem_b1_b_143 ), .B (n_5280), .S0 (n_5405), .Y(n_5281));
AOI22X1 g37317(.A0 (n_4729), .A1 (oc5_cfg_1015), .B0 (n_5591), .B1(n_4738), .Y (n_4741));
AOI22X1 g37316(.A0 (n_5272), .A1 (u13_intm_r_b10_b ), .B0 (n_5277),.B1 (crac_din_701), .Y (n_5279));
NAND2X1 g39071(.A (n_11804), .B (u8_mem_b0_b_111 ), .Y (n_3473));
INVX2 g40529(.A (wb_din_663), .Y (n_2804));
NAND2X1 g39076(.A (n_11798), .B (u8_mem_b0_b_104 ), .Y (n_11457));
NOR2X1 g41708(.A (n_705), .B (n_746), .Y (n_748));
NAND2X1 g39077(.A (u3_mem_b1_b_78 ), .B (n_3316), .Y (n_3469));
INVX4 g41707(.A (n_748), .Y (n_4961));
INVX4 g41706(.A (n_4961), .Y (n_1363));
NAND2X1 g39075(.A (u6_mem_b1_b ), .B (n_12169), .Y (n_11752));
INVX2 g45472(.A (n_12149), .Y (n_10787));
MX2X1 g40423(.A (crac_din_697), .B (in_slt_836), .S0 (n_1036), .Y(n_1196));
INVX2 g35032(.A (o3_we), .Y (n_8141));
INVX1 g35036(.A (n_7414), .Y (n_9333));
INVX1 g35037(.A (n_7414), .Y (n_9346));
INVX1 g35039(.A (n_7414), .Y (n_9336));
MX2X1 g36046(.A (n_6017), .B (n_6000), .S0 (n_6594), .Y (n_6001));
MX2X1 g36047(.A (n_6896), .B (n_6895), .S0 (n_6908), .Y (n_6897));
MX2X1 g36044(.A (n_6563), .B (n_6562), .S0 (n_6594), .Y (n_6564));
MX2X1 g36045(.A (n_6003), .B (n_6002), .S0 (n_6594), .Y (n_6004));
MX2X1 g36043(.A (n_6566), .B (n_6565), .S0 (n_6594), .Y (n_6567));
MX2X1 g36040(.A (n_6576), .B (n_6575), .S0 (n_6594), .Y (n_6577));
MX2X1 g36041(.A (n_6573), .B (n_6572), .S0 (n_6594), .Y (n_6574));
AOI21X1 g37768(.A0 (n_6426), .A1 (n_1831), .B0 (n_1005), .Y (n_1667));
INVX1 g42053(.A (u9_rp_b0_b ), .Y (n_121));
INVX1 g42050(.A (u9_mem_b1_b_140 ), .Y (n_1737));
INVX1 g42051(.A (u9_mem_b1_b_122 ), .Y (n_6876));
INVX1 g42059(.A (u11_mem_b3_b_60 ), .Y (n_6441));
NAND2X1 g37764(.A (n_3538), .B (n_2983), .Y (n_12850));
AOI22X1 g37765(.A0 (n_2502), .A1 (n_6854), .B0 (n_6876), .B1(n_1859), .Y (n_1669));
AOI22X1 g37766(.A0 (n_1756), .A1 (n_6370), .B0 (n_6517), .B1(n_1643), .Y (n_1668));
AOI21X1 g35960(.A0 (n_6972), .A1 (n_8528), .B0 (n_5784), .Y (n_6966));
AOI21X1 g35961(.A0 (n_6972), .A1 (n_8526), .B0 (n_5783), .Y (n_6965));
AOI21X1 g35962(.A0 (n_6972), .A1 (oc0_cfg_969), .B0 (n_5782), .Y(n_6964));
AOI21X1 g35963(.A0 (n_6972), .A1 (oc0_cfg_970), .B0 (n_5781), .Y(n_6963));
AOI21X1 g35964(.A0 (n_6972), .A1 (n_991), .B0 (n_5780), .Y (n_6962));
AOI21X1 g35965(.A0 (n_6972), .A1 (oc1_cfg_974), .B0 (n_5779), .Y(n_6961));
AOI21X1 g35966(.A0 (n_6972), .A1 (n_8567), .B0 (n_5761), .Y (n_6960));
AOI21X1 g35967(.A0 (n_6972), .A1 (oc1_cfg_975), .B0 (n_5786), .Y(n_6959));
AOI21X1 g35968(.A0 (n_6972), .A1 (oc1_cfg_979), .B0 (n_5777), .Y(n_6958));
MX2X1 g35969(.A (n_6037), .B (n_6017), .S0 (n_5407), .Y (n_6038));
NAND2X1 g39207(.A (u8_mem_b1_b_71 ), .B (n_12301), .Y (n_3374));
NOR2X1 g39201(.A (u10_mem_b1_b_133 ), .B (n_2364), .Y (n_2346));
NAND2X1 g39200(.A (u3_mem_b2_b_31 ), .B (n_12619), .Y (n_3383));
NOR2X1 g39202(.A (n_4961), .B (n_2765), .Y (n_3381));
NAND2X1 g39848(.A (n_2325), .B (in_slt_455), .Y (n_2238));
NAND2X1 g39843(.A (u3_mem_b1_b_67 ), .B (n_3316), .Y (n_2927));
OAI21X1 g35895(.A0 (n_5550), .A1 (n_7187), .B0 (n_6232), .Y (n_7094));
NOR2X1 g40299(.A (n_2025), .B (n_2702), .Y (n_1977));
NOR2X1 g39841(.A (n_3117), .B (n_2716), .Y (n_2929));
NOR2X1 g39840(.A (n_2748), .B (n_1488), .Y (n_1466));
NAND2X1 g39847(.A (n_2344), .B (in_slt_426), .Y (n_2239));
NAND2X1 g39846(.A (n_12369), .B (u6_mem_b0_b_99 ), .Y (n_2925));
NAND2X1 g34783(.A (u7_mem_b3_b_132 ), .B (n_7651), .Y (n_7650));
NAND2X1 g34782(.A (u7_mem_b3_b_131 ), .B (n_7651), .Y (n_7652));
NAND2X1 g34781(.A (u7_mem_b3_b ), .B (n_7651), .Y (n_7653));
NAND2X1 g34780(.A (u7_mem_b2_b_37 ), .B (n_7651), .Y (n_7654));
NAND2X1 g34787(.A (u7_mem_b3_b_136 ), .B (n_7651), .Y (n_7646));
NAND2X1 g34786(.A (u7_mem_b3_b_135 ), .B (n_7651), .Y (n_7647));
NAND2X1 g34785(.A (u7_mem_b3_b_134 ), .B (n_7651), .Y (n_7648));
NAND2X1 g34784(.A (u7_mem_b3_b_133 ), .B (n_7651), .Y (n_7649));
NAND2X1 g34789(.A (u7_mem_b3_b_138 ), .B (n_7651), .Y (n_7644));
NAND2X1 g34788(.A (u7_mem_b3_b_137 ), .B (n_7651), .Y (n_7645));
INVX1 g42701(.A (u10_mem_b0_b_164 ), .Y (n_6390));
NAND2X1 g34569(.A (u5_mem_b3_b_143 ), .B (n_7870), .Y (n_7857));
NAND2X1 g34568(.A (u5_mem_b3_b_142 ), .B (n_7870), .Y (n_7858));
NAND2X1 g34567(.A (u5_mem_b3_b_141 ), .B (n_7870), .Y (n_7859));
NAND2X1 g34566(.A (u5_mem_b3_b_122 ), .B (n_7870), .Y (n_7860));
NAND2X1 g34565(.A (u5_mem_b3_b_140 ), .B (n_7870), .Y (n_7861));
NAND2X1 g34564(.A (u5_mem_b3_b_139 ), .B (n_7870), .Y (n_7862));
NAND2X1 g34563(.A (u5_mem_b3_b_138 ), .B (n_7870), .Y (n_7863));
NAND2X1 g34562(.A (u5_mem_b3_b_137 ), .B (n_7870), .Y (n_7864));
NAND2X1 g34561(.A (u5_mem_b3_b_136 ), .B (n_7870), .Y (n_7865));
NAND2X1 g34560(.A (u5_mem_b3_b_135 ), .B (n_7870), .Y (n_7866));
INVX2 g43097(.A (u9_wp_b1_b ), .Y (n_689));
INVX1 g43096(.A (n_689), .Y (n_4074));
INVX1 g43090(.A (u10_mem_b2_b ), .Y (n_5998));
INVX1 g43093(.A (oc2_int_set_711), .Y (n_665));
INVX1 g45600(.A (n_12261), .Y (n_12262));
INVX2 g45602(.A (n_12269), .Y (n_12265));
NOR2X1 g41764(.A (n_715), .B (n_294), .Y (n_753));
INVX4 g40675(.A (wb_din_670), .Y (n_2691));
NAND2X1 g38958(.A (u7_mem_b3_b_137 ), .B (n_1546), .Y (n_1395));
NOR2X1 g40290(.A (n_941), .B (n_2741), .Y (n_1984));
NAND2X1 g38959(.A (u3_mem_b3_b_132 ), .B (n_2463), .Y (n_2397));
NAND2X1 g39812(.A (u7_mem_b2_b_31 ), .B (n_12645), .Y (n_2945));
INVX1 g42218(.A (u9_mem_b0_b_155 ), .Y (n_6849));
INVX1 g42874(.A (u10_mem_b3_b_71 ), .Y (n_6585));
INVX1 g42876(.A (u10_mem_b2_b_101 ), .Y (n_6662));
INVX1 g42877(.A (u15_crac_rd), .Y (n_36));
NAND2X1 g37148(.A (n_3938), .B (n_3348), .Y (n_6539));
NAND2X1 g37149(.A (n_2561), .B (n_4220), .Y (n_6618));
NAND2X1 g37144(.A (n_4626), .B (n_2354), .Y (n_6883));
NAND2X1 g37145(.A (n_3933), .B (n_3466), .Y (n_6582));
NAND2X1 g37146(.A (n_3934), .B (n_3081), .Y (n_6637));
NAND2X1 g37147(.A (n_3937), .B (n_3223), .Y (n_6533));
NAND2X1 g37141(.A (n_4619), .B (n_3373), .Y (n_6916));
NAND2X1 g37142(.A (n_3932), .B (n_1925), .Y (n_6560));
NAND2X1 g37143(.A (n_4625), .B (n_2259), .Y (n_6952));
NAND2X1 g36549(.A (n_12411), .B (n_6773), .Y (n_6771));
NAND2X1 g36548(.A (n_6147), .B (n_6773), .Y (n_6206));
NOR2X1 g36542(.A (i6_status), .B (n_11762), .Y (n_5434));
NAND2X1 g36541(.A (n_6209), .B (n_6773), .Y (n_6210));
NOR2X1 g36540(.A (i4_status), .B (n_11597), .Y (n_5594));
NAND2X1 g36547(.A (n_6773), .B (n_6769), .Y (n_6772));
NAND2X1 g36546(.A (n_6773), .B (n_6763), .Y (n_6774));
NAND4X1 g36545(.A (n_1014), .B (n_680), .C (u26_ps_cnt_b5_b ), .D(u26_ps_cnt_b4_b ), .Y (n_5632));
NAND2X1 g36544(.A (n_6207), .B (n_6773), .Y (n_6208));
INVX1 g42919(.A (n_431), .Y (n_4683));
INVX1 g42912(.A (u10_mem_b1_b_122 ), .Y (n_6542));
INVX1 g42911(.A (u9_mem_b3_b_80 ), .Y (n_5333));
INVX1 g42910(.A (u11_mem_b3_b_69 ), .Y (n_6424));
INVX1 g42916(.A (u10_mem_b2_b_90 ), .Y (n_6633));
INVX1 g42915(.A (u9_mem_b3_b_66 ), .Y (n_6620));
INVX1 g42914(.A (u9_mem_b3_b_68 ), .Y (n_6614));
INVX2 g45605(.A (n_12273), .Y (n_12269));
NOR2X1 g40734(.A (u10_rp_b1_b ), .B (n_403), .Y (n_940));
NOR2X1 g40988(.A (n_808), .B (n_4711), .Y (n_6201));
NOR2X1 g40209(.A (n_2171), .B (n_2792), .Y (n_2040));
INVX1 g45608(.A (n_12281), .Y (n_12274));
NAND2X1 g41242(.A (n_5), .B (n_487), .Y (n_603));
NOR2X1 g41243(.A (u13_ints_r_b16_b ), .B (n_463), .Y (n_696));
NOR2X1 g41240(.A (u9_rp_b0_b ), .B (n_4074), .Y (n_1054));
INVX2 g41241(.A (n_603), .Y (n_1756));
INVX1 g41647(.A (n_2468), .Y (n_1367));
OAI21X1 g31018(.A0 (n_5419), .A1 (n_10679), .B0 (n_9993), .Y(n_10678));
OAI21X1 g31019(.A0 (n_5428), .A1 (n_10820), .B0 (n_10393), .Y(n_10899));
INVX1 g42456(.A (u9_mem_b2_b_111 ), .Y (n_347));
OAI21X1 g31010(.A0 (n_5515), .A1 (n_10679), .B0 (n_10006), .Y(n_10690));
OAI21X1 g31011(.A0 (n_5513), .A1 (n_10679), .B0 (n_10005), .Y(n_10688));
OAI21X1 g31012(.A0 (n_5360), .A1 (n_10679), .B0 (n_10004), .Y(n_10686));
OAI21X1 g31013(.A0 (n_5358), .A1 (n_10450), .B0 (n_10003), .Y(n_10685));
OAI21X1 g31014(.A0 (n_5353), .A1 (n_10450), .B0 (n_10002), .Y(n_10684));
OAI21X1 g31015(.A0 (n_5511), .A1 (n_10450), .B0 (n_10001), .Y(n_10682));
OAI21X1 g31016(.A0 (n_5507), .A1 (n_10450), .B0 (n_10000), .Y(n_10681));
OAI21X1 g31017(.A0 (n_5505), .A1 (n_10679), .B0 (n_9999), .Y(n_10680));
NAND4X1 g33349(.A (n_5616), .B (n_1926), .C (n_7493), .D (n_1444), .Y(n_9449));
INVX4 g33342(.A (n_12503), .Y (n_10617));
NOR2X1 g41060(.A (n_621), .B (wb_addr_i_b3_b), .Y (n_6044));
OR2X1 g41066(.A (n_590), .B (oc5_cfg_1016), .Y (n_6981));
NAND2X1 g40984(.A (n_145), .B (n_765), .Y (n_929));
INVX2 g41064(.A (n_1038), .Y (n_7063));
INVX1 g41065(.A (n_6981), .Y (n_1038));
MX2X1 g31274(.A (n_6850), .B (n_6849), .S0 (n_10250), .Y (n_10145));
MX2X1 g31275(.A (n_6848), .B (n_6847), .S0 (n_10250), .Y (n_10143));
MX2X1 g31276(.A (n_6395), .B (n_6394), .S0 (n_10250), .Y (n_10142));
MX2X1 g31277(.A (n_6846), .B (n_6845), .S0 (n_10235), .Y (n_10141));
MX2X1 g31270(.A (n_6858), .B (n_6857), .S0 (n_10267), .Y (n_10148));
MX2X1 g31271(.A (n_6855), .B (n_6854), .S0 (n_10267), .Y (n_10147));
XOR2X1 g31272(.A (n_634), .B (n_9907), .Y (n_10822));
MX2X1 g31273(.A (n_6853), .B (n_6852), .S0 (n_10267), .Y (n_10146));
OAI21X1 g31278(.A0 (n_10992), .A1 (u4_rp_b0_b ), .B0 (n_9843), .Y(n_10140));
OAI21X1 g31279(.A0 (n_10985), .A1 (n_5772), .B0 (n_9842), .Y(n_10139));
INVX2 g42454(.A (u10_rp_b0_b ), .Y (n_403));
OAI21X1 g33954(.A0 (n_4861), .A1 (n_8911), .B0 (n_7947), .Y (n_8874));
OAI21X1 g33518(.A0 (n_4461), .A1 (n_8333), .B0 (n_8041), .Y (n_8329));
NAND2X1 g34673(.A (u6_mem_b3_b_138 ), .B (n_7758), .Y (n_7751));
INVX2 g40985(.A (n_6201), .Y (n_7088));
OAI21X1 g33952(.A0 (n_4500), .A1 (n_8898), .B0 (n_8076), .Y (n_8876));
NOR2X1 g40195(.A (n_2133), .B (n_2790), .Y (n_2049));
NAND2X1 g34671(.A (u6_mem_b3_b_136 ), .B (n_7758), .Y (n_7753));
NAND2X1 g36364(.A (n_5815), .B (n_2567), .Y (n_5916));
INVX1 g40719(.A (n_1176), .Y (n_2093));
NAND2X1 g38964(.A (u7_mem_b3_b_138 ), .B (n_1546), .Y (n_1376));
NAND2X1 g34248(.A (u8_mem_b3_b_140 ), .B (n_7976), .Y (n_8154));
OAI21X1 g33569(.A0 (n_4408), .A1 (n_8333), .B0 (n_7988), .Y (n_8267));
OAI21X1 g33959(.A0 (n_4396), .A1 (n_8868), .B0 (n_7571), .Y (n_8867));
INVX2 g41351(.A (n_1134), .Y (n_6908));
OAI21X1 g33958(.A0 (n_4291), .A1 (n_8868), .B0 (n_7616), .Y (n_8869));
INVX1 g40689(.A (n_1180), .Y (n_2118));
INVX1 g40688(.A (n_1180), .Y (n_2057));
INVX1 g41353(.A (n_1134), .Y (n_1063));
AND2X1 g41354(.A (u9_wp_b1_b ), .B (u9_wp_b2_b ), .Y (n_1134));
INVX4 g40682(.A (wb_din_682), .Y (n_2792));
BUFX3 g40685(.A (n_933), .Y (n_4387));
BUFX3 g40684(.A (n_933), .Y (n_4502));
INVX1 g40687(.A (n_1180), .Y (n_2008));
OAI21X1 g33787(.A0 (n_5060), .A1 (n_9087), .B0 (n_7740), .Y (n_9088));
OAI21X1 g33562(.A0 (n_4417), .A1 (n_9336), .B0 (n_7995), .Y (n_8274));
NAND2X1 g36369(.A (n_5694), .B (n_12634), .Y (n_6300));
CLKBUFX1 g41357(.A (n_1064), .Y (n_5645));
NAND2X1 g34240(.A (u8_mem_b3_b_132 ), .B (n_7976), .Y (n_8165));
CLKBUFX2 g40922(.A (n_932), .Y (n_5409));
OAI21X1 g33561(.A0 (n_4418), .A1 (n_8333), .B0 (n_7996), .Y (n_8275));
OAI21X1 g33566(.A0 (n_4411), .A1 (n_8333), .B0 (n_7991), .Y (n_8270));
OAI21X1 g33567(.A0 (n_4410), .A1 (n_8333), .B0 (n_7990), .Y (n_8269));
NAND3X1 g30053(.A (n_9698), .B (n_9523), .C (n_9655), .Y (n_9848));
NAND3X1 g30052(.A (n_9767), .B (n_9600), .C (n_9658), .Y (n_10091));
NAND3X1 g30051(.A (n_9700), .B (n_9524), .C (n_9613), .Y (n_9849));
AOI21X1 g35570(.A0 (n_6326), .A1 (n_6129), .B0 (n_7324), .Y (n_7275));
OAI21X1 g30057(.A0 (n_9504), .A1 (n_9589), .B0 (n_9755), .Y(n_10089));
AOI21X1 g35575(.A0 (n_6833), .A1 (n_6126), .B0 (n_7324), .Y (n_7325));
NAND3X1 g30054(.A (n_9696), .B (n_9522), .C (n_9652), .Y (n_9847));
NOR2X1 g39018(.A (n_3089), .B (n_2686), .Y (n_3512));
NOR2X1 g39019(.A (n_3486), .B (n_2732), .Y (n_3511));
AOI21X1 g35579(.A0 (n_11539), .A1 (n_11540), .B0 (n_12145), .Y(n_7320));
OAI21X1 g30058(.A0 (n_9561), .A1 (n_9645), .B0 (n_9837), .Y(n_10400));
NAND4X1 g36848(.A (n_4192), .B (n_1491), .C (n_2314), .D (n_4257), .Y(n_6807));
INVX1 g36849(.A (n_6800), .Y (n_6078));
NAND2X1 g36846(.A (n_1695), .B (n_3929), .Y (n_5393));
INVX1 g36847(.A (n_6807), .Y (n_6079));
INVX1 g36844(.A (n_6803), .Y (n_6080));
NAND4X1 g36845(.A (n_4195), .B (n_3108), .C (n_2277), .D (n_4259), .Y(n_6803));
NAND4X1 g36842(.A (n_4144), .B (n_2972), .C (n_2260), .D (n_4252), .Y(n_6797));
NAND4X1 g36843(.A (n_4147), .B (n_3393), .C (n_2348), .D (n_4260), .Y(n_6794));
INVX1 g36840(.A (n_6790), .Y (n_6081));
NAND4X1 g36841(.A (n_4243), .B (n_3517), .C (n_2350), .D (n_4261), .Y(n_6790));
INVX1 g34998(.A (n_7424), .Y (n_9022));
INVX1 g34999(.A (n_7424), .Y (n_8375));
INVX1 g34996(.A (n_7424), .Y (n_8372));
INVX1 g34997(.A (n_7424), .Y (n_8369));
INVX1 g34994(.A (n_7424), .Y (n_8380));
INVX1 g34995(.A (n_7424), .Y (n_8383));
INVX1 g34992(.A (n_7424), .Y (n_8387));
INVX1 g34993(.A (n_7424), .Y (n_8357));
INVX1 g37416(.A (n_3945), .Y (n_4679));
INVX1 g45604(.A (n_12269), .Y (n_12270));
XOR2X1 g37417(.A (u8_wp_b1_b ), .B (n_12278), .Y (n_1294));
AOI22X1 g37946(.A0 (n_2558), .A1 (n_5957), .B0 (n_5974), .B1(n_1839), .Y (n_2504));
NAND2X1 g37940(.A (n_2432), .B (n_3315), .Y (n_5194));
NAND2X1 g36418(.A (n_6165), .B (n_12115), .Y (n_6263));
AOI22X1 g37942(.A0 (u11_din_tmp_56), .A1 (n_4560), .B0 (n_4097), .B1(in_slt_457), .Y (n_4098));
NAND2X1 g37943(.A (n_1525), .B (n_4128), .Y (n_5452));
MX2X1 g36146(.A (n_6849), .B (n_6899), .S0 (n_6856), .Y (n_6850));
OAI21X1 g33500(.A0 (n_5126), .A1 (n_8387), .B0 (n_7834), .Y (n_8352));
OAI21X1 g33501(.A0 (n_4527), .A1 (n_8894), .B0 (n_7592), .Y (n_8351));
OAI21X1 g33502(.A0 (n_3872), .A1 (n_8464), .B0 (n_8147), .Y (n_8350));
OAI21X1 g33503(.A0 (n_4485), .A1 (n_8891), .B0 (n_7558), .Y (n_8349));
OAI21X1 g33504(.A0 (n_4960), .A1 (n_9022), .B0 (n_8086), .Y (n_8348));
OAI21X1 g33505(.A0 (n_4855), .A1 (n_8911), .B0 (n_7559), .Y (n_8347));
OAI21X1 g33506(.A0 (n_4345), .A1 (n_8393), .B0 (n_8066), .Y (n_8346));
OAI21X1 g33507(.A0 (n_4473), .A1 (n_8333), .B0 (n_8056), .Y (n_8345));
OAI21X1 g33508(.A0 (n_4381), .A1 (n_9349), .B0 (n_8055), .Y (n_8344));
OAI21X1 g33509(.A0 (n_4472), .A1 (n_8333), .B0 (n_8054), .Y (n_8343));
NAND2X1 g36410(.A (n_6839), .B (n_6838), .Y (n_5901));
INVX1 g41972(.A (u11_mem_b1_b_147 ), .Y (n_1591));
NAND2X1 g36413(.A (n_6264), .B (n_6201), .Y (n_6265));
MX2X1 g36140(.A (n_6864), .B (n_6952), .S0 (n_6856), .Y (n_6865));
NAND2X1 g37557(.A (n_5656), .B (n_4138), .Y (n_5239));
NAND2X1 g37556(.A (n_5645), .B (n_4111), .Y (n_5240));
NAND2X1 g37555(.A (n_5656), .B (n_4237), .Y (n_5241));
NAND2X1 g37554(.A (n_5656), .B (n_4205), .Y (n_5242));
NOR2X1 g37553(.A (n_4757), .B (n_5371), .Y (n_3949));
NOR2X1 g37552(.A (n_5296), .B (n_6649), .Y (n_4643));
NOR2X1 g37551(.A (n_4776), .B (n_5371), .Y (n_3950));
OAI21X1 g37550(.A0 (n_1205), .A1 (u5_rp_b3_b ), .B0 (n_4644), .Y(n_4645));
NAND2X1 g37559(.A (n_5645), .B (n_2994), .Y (n_4642));
NAND2X1 g37558(.A (n_5656), .B (n_4202), .Y (n_5238));
OAI21X1 g33647(.A0 (n_4368), .A1 (n_9212), .B0 (n_7893), .Y (n_9261));
OAI21X1 g33646(.A0 (n_4276), .A1 (n_9288), .B0 (n_7894), .Y (n_9262));
OAI21X1 g33645(.A0 (n_4369), .A1 (n_9307), .B0 (n_7895), .Y (n_9263));
OAI21X1 g33644(.A0 (n_4371), .A1 (n_9264), .B0 (n_7896), .Y (n_9265));
OAI21X1 g33643(.A0 (n_4372), .A1 (n_9307), .B0 (n_7897), .Y (n_9266));
OAI21X1 g33642(.A0 (n_4373), .A1 (n_9290), .B0 (n_7898), .Y (n_9267));
OAI21X1 g33641(.A0 (n_4374), .A1 (n_9307), .B0 (n_7899), .Y (n_9268));
OAI21X1 g33640(.A0 (n_4542), .A1 (n_9288), .B0 (n_7900), .Y (n_9269));
NAND4X1 g37081(.A (n_12827), .B (n_12828), .C (n_2246), .D (n_3539),.Y (n_6180));
INVX1 g37080(.A (n_6180), .Y (n_5678));
NAND4X1 g37083(.A (n_3375), .B (n_3199), .C (n_3119), .D (n_1508), .Y(n_6144));
INVX1 g37082(.A (n_6144), .Y (n_5677));
NAND4X1 g37085(.A (n_11467), .B (n_11468), .C (n_2245), .D (n_2395),.Y (n_5803));
INVX1 g37084(.A (n_5803), .Y (n_5536));
OAI21X1 g33649(.A0 (n_4365), .A1 (n_9288), .B0 (n_7891), .Y (n_9258));
OAI21X1 g33648(.A0 (n_4367), .A1 (n_9290), .B0 (n_7892), .Y (n_9259));
NAND2X1 g39628(.A (n_12204), .B (u6_mem_b0_b_109 ), .Y (n_12817));
INVX4 g40536(.A (wb_din_662), .Y (n_2782));
NAND2X1 g38962(.A (u8_mem_b3_b_135 ), .B (n_2468), .Y (n_1892));
NOR2X1 g34702(.A (o9_status_1012), .B (n_12585), .Y (n_9481));
INVX1 g42381(.A (n_9833), .Y (n_10994));
AOI22X1 g37333(.A0 (n_5272), .A1 (u13_intm_r_b22_b ), .B0(u13_ints_r_b22_b ), .B1 (n_4726), .Y (n_4722));
OAI21X1 g33481(.A0 (n_5132), .A1 (n_8372), .B0 (n_8090), .Y (n_8374));
INVX1 g37331(.A (n_3989), .Y (n_4723));
NAND2X1 g37882(.A (n_4143), .B (n_3041), .Y (n_5197));
AOI22X1 g37337(.A0 (n_5272), .A1 (u13_intm_r_b24_b ), .B0 (n_6972),.B1 (n_1873), .Y (n_4719));
AOI21X1 g38500(.A0 (u7_mem_b2_b_54 ), .A1 (n_4509), .B0 (n_1977), .Y(n_4311));
INVX1 g37335(.A (n_3986), .Y (n_4720));
NAND2X1 g34452(.A (u4_mem_b3_b_142 ), .B (n_7984), .Y (n_7969));
AOI22X1 g37889(.A0 (u11_din_tmp_54), .A1 (n_4560), .B0 (n_4097), .B1(in_slt_455), .Y (n_3902));
AOI22X1 g37888(.A0 (n_1756), .A1 (n_6372), .B0 (n_6519), .B1(n_1643), .Y (n_1837));
AOI22X1 g37339(.A0 (n_5272), .A1 (u13_intm_r_b26_b ), .B0 (n_6972),.B1 (oc3_cfg_995), .Y (n_5274));
AOI22X1 g37338(.A0 (n_5272), .A1 (u13_intm_r_b25_b ), .B0 (n_6972),.B1 (oc3_cfg_994), .Y (n_4718));
AOI21X1 g38509(.A0 (u7_mem_b2_b_37 ), .A1 (n_4540), .B0 (n_2019), .Y(n_4303));
OAI21X1 g33483(.A0 (n_5093), .A1 (n_8369), .B0 (n_8087), .Y (n_8371));
INVX2 g41139(.A (n_1411), .Y (n_3423));
AOI21X1 g34906(.A0 (n_4102), .A1 (n_2513), .B0 (n_2606), .Y (n_5634));
MX2X1 g38737(.A (u3_mem_b0_b_106 ), .B (wb_din_676), .S0 (n_3807), .Y(n_3603));
NAND2X1 g34457(.A (u4_mem_b3_b_147 ), .B (n_7984), .Y (n_7964));
OAI21X1 g33484(.A0 (n_5131), .A1 (n_8369), .B0 (n_8061), .Y (n_8370));
MX2X1 g36091(.A (n_6487), .B (n_6486), .S0 (n_6502), .Y (n_6488));
OAI21X1 g33487(.A0 (n_5123), .A1 (n_8369), .B0 (n_8084), .Y (n_8366));
NAND2X1 g34454(.A (u4_mem_b3_b_144 ), .B (n_7984), .Y (n_7967));
INVX2 g39672(.A (n_1216), .Y (n_5277));
OAI21X1 g36684(.A0 (n_5171), .A1 (n_4580), .B0 (n_6152), .Y (n_5759));
OAI21X1 g36680(.A0 (n_5461), .A1 (n_5205), .B0 (n_6118), .Y (n_6106));
OAI21X1 g36681(.A0 (n_4610), .A1 (n_5197), .B0 (n_784), .Y (n_6105));
OAI21X1 g36682(.A0 (n_12060), .A1 (n_12061), .B0 (n_784), .Y(n_6104));
OAI21X1 g36683(.A0 (n_5170), .A1 (n_5168), .B0 (n_634), .Y (n_5760));
OAI21X1 g36688(.A0 (n_4574), .A1 (n_5172), .B0 (n_6152), .Y (n_5758));
NAND2X1 g45794(.A (n_12641), .B (u7_mem_b2_b_32 ), .Y (n_12513));
NAND4X1 g45790(.A (n_12506), .B (n_12507), .C (n_12508), .D(n_12513), .Y (n_12514));
NAND2X1 g45791(.A (n_4130), .B (u7_mem_b1_b_63 ), .Y (n_12506));
NAND2X1 g45793(.A (n_1538), .B (u7_mem_b3_b_125 ), .Y (n_12508));
NAND2X1 g45798(.A (n_438), .B (n_12330), .Y (n_12509));
AOI21X1 g30736(.A0 (n_9768), .A1 (n_9660), .B0 (n_9648), .Y (n_9769));
AOI21X1 g30737(.A0 (n_9699), .A1 (n_9612), .B0 (n_9590), .Y (n_9700));
AOI21X1 g30734(.A0 (n_7519), .A1 (n_9444), .B0 (n_9526), .Y(n_11504));
AOI21X1 g30735(.A0 (n_9701), .A1 (n_9615), .B0 (n_9592), .Y (n_9702));
AOI21X1 g30732(.A0 (n_7448), .A1 (n_8847), .B0 (n_9474), .Y(n_11672));
AOI21X1 g30733(.A0 (n_7446), .A1 (n_8843), .B0 (n_9473), .Y(n_11673));
OR2X1 g30730(.A (n_10403), .B (n_11131), .Y (n_11510));
OR2X1 g30731(.A (n_10402), .B (n_11126), .Y (n_11508));
AOI21X1 g30738(.A0 (n_9766), .A1 (n_9657), .B0 (n_9646), .Y (n_9767));
AOI21X1 g30739(.A0 (n_9697), .A1 (n_9654), .B0 (n_9588), .Y (n_9698));
INVX4 g41476(.A (n_4996), .Y (n_1388));
NOR2X1 g40274(.A (n_2038), .B (n_2681), .Y (n_1995));
INVX1 g35015(.A (n_7424), .Y (n_8393));
INVX1 g35017(.A (n_7424), .Y (n_8440));
NOR2X1 g41479(.A (wb_addr_i_b2_b), .B (wb_addr_i_b3_b), .Y (n_996));
NOR2X1 g41478(.A (n_734), .B (n_710), .Y (n_615));
INVX2 g35012(.A (n_7424), .Y (n_8911));
MX2X1 g36060(.A (n_6542), .B (n_6573), .S0 (n_832), .Y (n_6543));
MX2X1 g36061(.A (n_6540), .B (n_6539), .S0 (n_4783), .Y (n_6541));
MX2X1 g36062(.A (n_6537), .B (n_6560), .S0 (n_5730), .Y (n_6538));
MX2X1 g36063(.A (n_508), .B (n_6589), .S0 (n_6475), .Y (n_6536));
MX2X1 g36064(.A (n_6534), .B (n_6533), .S0 (n_4783), .Y (n_6535));
MX2X1 g36066(.A (n_6879), .B (n_6916), .S0 (n_4783), .Y (n_6880));
MX2X1 g36067(.A (n_6876), .B (n_6896), .S0 (n_969), .Y (n_6877));
MX2X1 g36068(.A (n_6530), .B (n_6547), .S0 (n_5312), .Y (n_6531));
MX2X1 g36069(.A (n_6528), .B (n_6582), .S0 (n_4783), .Y (n_6529));
NOR2X1 g40017(.A (n_2832), .B (n_2818), .Y (n_2819));
INVX1 g42079(.A (u9_mem_b2_b_95 ), .Y (n_6628));
INVX1 g42074(.A (u11_mem_b0_b_176 ), .Y (n_1600));
INVX1 g42076(.A (u11_mem_b2_b_111 ), .Y (n_275));
INVX1 g42071(.A (u14_n_133), .Y (n_1308));
NAND3X1 g45747(.A (n_12535), .B (n_6316), .C (n_12111), .Y (n_12459));
NAND2X1 g34629(.A (u6_mem_b1_b_66 ), .B (n_7758), .Y (n_7796));
NOR2X1 g35337(.A (n_6046), .B (u2_bit_clk_e), .Y (n_7033));
OAI21X1 g35908(.A0 (n_5671), .A1 (n_7088), .B0 (n_6234), .Y (n_7087));
OAI21X1 g35909(.A0 (n_5691), .A1 (n_7088), .B0 (n_6210), .Y (n_7085));
NAND2X1 g39676(.A (u5_mem_b1_b_76 ), .B (n_3236), .Y (n_11482));
OAI21X1 g35902(.A0 (n_5547), .A1 (n_7187), .B0 (n_5834), .Y (n_6990));
OAI21X1 g35903(.A0 (n_5555), .A1 (n_7187), .B0 (n_5856), .Y (n_6989));
OAI21X1 g35900(.A0 (n_5702), .A1 (n_7187), .B0 (n_5838), .Y (n_7092));
OAI21X1 g35901(.A0 (n_5548), .A1 (n_7187), .B0 (n_5836), .Y (n_6991));
OAI21X1 g35906(.A0 (n_5545), .A1 (n_7088), .B0 (n_6215), .Y (n_7090));
OAI21X1 g35907(.A0 (n_5692), .A1 (n_7088), .B0 (n_6212), .Y (n_7089));
OAI21X1 g35904(.A0 (n_5553), .A1 (n_7187), .B0 (n_6780), .Y (n_7183));
OAI21X1 g35905(.A0 (n_5693), .A1 (n_7088), .B0 (n_6217), .Y (n_7091));
INVX1 g41644(.A (n_12603), .Y (n_7267));
NOR2X1 g35336(.A (n_5614), .B (u2_bit_clk_e), .Y (n_6733));
NOR2X1 g40277(.A (n_2477), .B (n_2729), .Y (n_1992));
INVX1 g42593(.A (u10_mem_b2_b_115 ), .Y (n_2545));
NAND2X1 g34769(.A (u7_mem_b2_b_56 ), .B (n_7651), .Y (n_7665));
NAND2X1 g34768(.A (u7_mem_b2_b_55 ), .B (n_7651), .Y (n_7666));
NAND2X1 g34765(.A (u7_mem_b2_b_52 ), .B (n_7651), .Y (n_7669));
NAND2X1 g34764(.A (u7_mem_b2_b_51 ), .B (n_7651), .Y (n_7670));
NAND2X1 g34767(.A (u7_mem_b2_b_54 ), .B (n_7651), .Y (n_7667));
NAND2X1 g34766(.A (u7_mem_b2_b_53 ), .B (n_7651), .Y (n_7668));
NAND2X1 g34760(.A (u7_mem_b2_b_47 ), .B (n_7651), .Y (n_7674));
NAND2X1 g34763(.A (u7_mem_b2_b_50 ), .B (n_7651), .Y (n_7671));
NAND2X1 g34762(.A (u7_mem_b2_b_49 ), .B (n_7651), .Y (n_7672));
NOR2X1 g39227(.A (u10_mem_b1_b_135 ), .B (n_2364), .Y (n_2365));
NAND2X1 g39226(.A (u8_mem_b1_b_64 ), .B (n_12291), .Y (n_3355));
NAND2X1 g39225(.A (u6_mem_b1_b_90 ), .B (n_12169), .Y (n_4212));
NAND2X1 g39224(.A (n_2344), .B (in_slt_433), .Y (n_2345));
NAND2X1 g39223(.A (u7_mem_b1_b_85 ), .B (n_4225), .Y (n_4214));
NOR2X1 g39222(.A (n_3332), .B (n_2735), .Y (n_3357));
NOR2X1 g39221(.A (n_3089), .B (n_2767), .Y (n_3358));
NAND2X1 g39220(.A (u8_mem_b2_b_42 ), .B (n_2362), .Y (n_2128));
INVX1 g42598(.A (u11_mem_b1_b_141 ), .Y (n_1619));
INVX1 g41687(.A (n_1107), .Y (n_1364));
NOR2X1 g39229(.A (n_3117), .B (n_2782), .Y (n_3353));
INVX1 g41830(.A (u11_mem_b1_b_140 ), .Y (n_1754));
INVX1 g41811(.A (u11_mem_b0_b_164 ), .Y (n_6360));
INVX1 g41810(.A (u10_mem_b3_b_82 ), .Y (n_5359));
INVX1 g40840(.A (n_1167), .Y (n_2041));
NAND2X1 g34509(.A (u5_mem_b1_b_86 ), .B (n_7870), .Y (n_7919));
NAND2X1 g34508(.A (u5_mem_b1_b_85 ), .B (n_7870), .Y (n_7920));
INVX4 g40659(.A (wb_din_675), .Y (n_2741));
AOI21X1 g38521(.A0 (u7_mem_b3_b_150 ), .A1 (n_4961), .B0 (n_3417), .Y(n_4880));
INVX1 g35332(.A (n_7536), .Y (n_8679));
NAND2X1 g34501(.A (u5_mem_b1_b_60 ), .B (n_7870), .Y (n_7929));
NAND2X1 g34500(.A (u5_mem_b1_b_78 ), .B (n_7870), .Y (n_7930));
NAND2X1 g34503(.A (u5_mem_b1_b_80 ), .B (n_7870), .Y (n_7925));
NAND2X1 g34505(.A (u5_mem_b1_b_82 ), .B (n_7870), .Y (n_7923));
NAND2X1 g34504(.A (u5_mem_b1_b_81 ), .B (n_7870), .Y (n_7924));
NAND2X1 g34507(.A (u5_mem_b1_b_84 ), .B (n_7870), .Y (n_7921));
NAND2X1 g34506(.A (u5_mem_b1_b_83 ), .B (n_7870), .Y (n_7922));
OAI21X1 g33470(.A0 (n_4859), .A1 (n_8387), .B0 (n_8104), .Y (n_8389));
OAI21X1 g45740(.A0 (n_12454), .A1 (n_12460), .B0 (n_10481), .Y(n_12464));
NAND2X1 g39736(.A (u9_din_tmp_50), .B (n_2368), .Y (n_2255));
NOR2X1 g40845(.A (n_8550), .B (n_503), .Y (n_9699));
NAND2X1 g38818(.A (u6_mem_b3_b_130 ), .B (n_12622), .Y (n_1861));
NOR2X1 g39731(.A (n_5102), .B (n_2772), .Y (n_2992));
NAND2X1 g45884(.A (n_12825), .B (u3_mem_b0_b_102 ), .Y (n_12612));
NAND2X1 g45885(.A (n_1517), .B (u3_mem_b3_b_133 ), .Y (n_12613));
NOR2X1 g39836(.A (n_3117), .B (n_2681), .Y (n_2932));
OAI21X1 g33475(.A0 (n_4955), .A1 (n_8380), .B0 (n_8096), .Y (n_8382));
NAND4X1 g36827(.A (n_11656), .B (n_11657), .C (n_3248), .D (n_3547),.Y (n_6266));
INVX1 g42898(.A (u10_mem_b3_b_85 ), .Y (n_5510));
INVX1 g42899(.A (u10_mem_b2_b_105 ), .Y (n_1690));
INVX4 g42896(.A (u3_rp_b0_b ), .Y (n_6316));
NAND2X1 g39837(.A (n_12826), .B (u3_mem_b0_b_105 ), .Y (n_12834));
INVX4 g42895(.A (n_6316), .Y (n_634));
OAI21X1 g33871(.A0 (n_4303), .A1 (n_9055), .B0 (n_7654), .Y (n_8984));
NOR2X1 g40029(.A (n_2775), .B (n_2707), .Y (n_2814));
NOR2X1 g40028(.A (n_935), .B (n_2741), .Y (n_2188));
NOR2X1 g40024(.A (n_2831), .B (n_2182), .Y (n_2192));
NOR2X1 g40027(.A (n_1016), .B (n_2732), .Y (n_2815));
NOR2X1 g40026(.A (n_2189), .B (n_2786), .Y (n_2190));
NOR2X1 g40021(.A (n_2686), .B (n_1985), .Y (n_2196));
NOR2X1 g40020(.A (n_2773), .B (n_2829), .Y (n_2816));
NOR2X1 g40023(.A (n_2765), .B (n_2067), .Y (n_2193));
NOR2X1 g40022(.A (n_945), .B (n_2767), .Y (n_2195));
NAND2X1 g39834(.A (u8_mem_b1_b_62 ), .B (n_12301), .Y (n_11503));
INVX1 g36821(.A (n_6246), .Y (n_5728));
AOI22X1 g35506(.A0 (n_5630), .A1 (n_4088), .B0 (n_5629), .B1(n_4089), .Y (n_5614));
AOI21X1 g30027(.A0 (n_9555), .A1 (n_9699), .B0 (n_10089), .Y(n_10408));
XOR2X1 g35500(.A (n_6047), .B (n_4841), .Y (n_6048));
AND2X1 g30021(.A (n_11150), .B (n_9833), .Y (n_11164));
INVX1 g41897(.A (oc3_cfg_999), .Y (n_485));
INVX1 g41894(.A (u10_mem_b1_b_121 ), .Y (n_6415));
INVX1 g41892(.A (u9_mem_b0_b_160 ), .Y (n_6402));
INVX1 g41891(.A (u11_rp_b0_b ), .Y (n_487));
NAND2X1 g39891(.A (u8_mem_b2_b_34 ), .B (n_2362), .Y (n_2509));
MX2X1 g38741(.A (u8_mem_b0_b_106 ), .B (wb_din_676), .S0 (n_3826), .Y(n_3599));
NOR2X1 g41268(.A (u13_ints_r_b10_b ), .B (n_450), .Y (n_694));
INVX1 g41264(.A (n_695), .Y (n_914));
NAND2X1 g41265(.A (u11_wp_b1_b ), .B (u11_wp_b2_b ), .Y (n_695));
AND2X1 g41266(.A (n_598), .B (n_804), .Y (n_9650));
OAI21X1 g31072(.A0 (n_5501), .A1 (n_10820), .B0 (n_10350), .Y(n_10850));
OAI21X1 g31073(.A0 (n_5503), .A1 (n_10820), .B0 (n_10349), .Y(n_10849));
OAI21X1 g31070(.A0 (n_5497), .A1 (n_10820), .B0 (n_10352), .Y(n_10852));
OAI21X1 g31071(.A0 (n_5493), .A1 (n_10820), .B0 (n_10351), .Y(n_10851));
OAI21X1 g31076(.A0 (n_5509), .A1 (n_10880), .B0 (n_10346), .Y(n_10846));
OAI21X1 g31077(.A0 (n_5523), .A1 (n_10880), .B0 (n_10345), .Y(n_10845));
OAI21X1 g31074(.A0 (n_5499), .A1 (n_10820), .B0 (n_10348), .Y(n_10848));
OAI21X1 g31075(.A0 (n_5525), .A1 (n_10820), .B0 (n_10347), .Y(n_10847));
INVX1 g42791(.A (u11_wp_b2_b ), .Y (n_520));
INVX1 g42790(.A (n_520), .Y (n_853));
AOI21X1 g31078(.A0 (n_11893), .A1 (u8_rp_b3_b ), .B0 (n_9974), .Y(n_10663));
AOI21X1 g31079(.A0 (n_12339), .A1 (u3_rp_b3_b ), .B0 (n_9973), .Y(n_10661));
INVX1 g42794(.A (n_462), .Y (n_4710));
INVX1 g42797(.A (u10_mem_b3_b_67 ), .Y (n_6598));
INVX1 g42796(.A (ic0_cfg_1026), .Y (n_462));
AOI22X1 g37353(.A0 (n_4729), .A1 (n_4701), .B0 (n_5591), .B1(n_4699), .Y (n_4702));
INVX2 g41044(.A (n_1412), .Y (n_3239));
INVX4 g41045(.A (n_1035), .Y (n_1412));
INVX1 g41046(.A (n_3209), .Y (n_1908));
INVX1 g41047(.A (n_1412), .Y (n_3209));
INVX1 g33360(.A (n_9666), .Y (n_9703));
INVX1 g33361(.A (n_9567), .Y (n_9666));
NOR2X1 g33362(.A (n_11530), .B (n_8661), .Y (n_9567));
NAND4X1 g33363(.A (n_5622), .B (n_1929), .C (n_7490), .D (n_1447), .Y(n_9448));
INVX1 g33368(.A (n_9514), .Y (n_9690));
INVX2 g33369(.A (n_9447), .Y (n_9514));
AOI22X1 g40414(.A0 (u13_intm_r_b23_b ), .A1 (u13_ints_r_b23_b ), .B0(u13_intm_r_b24_b ), .B1 (u13_ints_r_b24_b ), .Y (n_729));
NAND2X1 g39894(.A (u3_mem_b2_b_59 ), .B (n_3330), .Y (n_2896));
NAND2X2 g40963(.A (n_798), .B (n_734), .Y (n_1082));
MX2X1 g38730(.A (u6_mem_b0_b_112 ), .B (wb_din_682), .S0 (n_3632), .Y(n_3611));
MX2X1 g31299(.A (n_5952), .B (n_5951), .S0 (n_10513), .Y (n_10447));
MX2X1 g31296(.A (n_5956), .B (n_5955), .S0 (n_10315), .Y (n_10131));
MX2X1 g31297(.A (n_5954), .B (n_5953), .S0 (n_10513), .Y (n_10448));
MX2X1 g31295(.A (n_6361), .B (n_6360), .S0 (n_9818), .Y (n_10813));
MX2X1 g31292(.A (n_5958), .B (n_5957), .S0 (n_10315), .Y (n_10132));
MX2X1 g31293(.A (n_6364), .B (n_6363), .S0 (n_9818), .Y (n_10814));
MX2X1 g31291(.A (n_6367), .B (n_6366), .S0 (n_9818), .Y (n_10817));
INVX1 g42123(.A (u10_mem_b2_b_89 ), .Y (n_6652));
NAND2X1 g39502(.A (in_slt_412), .B (n_2368), .Y (n_4772));
NAND2X1 g39500(.A (n_12840), .B (u4_mem_b0_b_104 ), .Y (n_11650));
AOI22X1 g40416(.A0 (u13_intm_r_b1_b ), .A1 (u13_ints_r_b1_b ), .B0(u13_intm_r_b3_b ), .B1 (u13_ints_r_b3_b ), .Y (n_792));
NAND2X1 g39896(.A (in_slt_405), .B (n_2368), .Y (n_4747));
INVX1 g39501(.A (n_4772), .Y (n_3138));
NAND2X1 g39506(.A (u3_mem_b1_b_61 ), .B (n_3316), .Y (n_3135));
NAND2X1 g39504(.A (in_slt_411), .B (n_2368), .Y (n_4743));
AOI22X1 g40417(.A0 (u13_intm_r_b19_b ), .A1 (u13_ints_r_b19_b ), .B0(u13_intm_r_b20_b ), .B1 (u13_ints_r_b20_b ), .Y (n_726));
NOR2X1 g39897(.A (n_2684), .B (n_1488), .Y (n_1462));
INVX1 g42449(.A (n_8565), .Y (n_693));
INVX1 g43042(.A (n_422), .Y (n_1873));
INVX1 g42241(.A (u11_mem_b2_b_103 ), .Y (n_5994));
INVX1 g42240(.A (u10_mem_b1_b_126 ), .Y (n_5966));
INVX1 g42531(.A (n_838), .Y (n_2574));
INVX1 g42246(.A (u9_mem_b2_b_98 ), .Y (n_6644));
INVX2 g42533(.A (wb_addr_i_b2_b), .Y (n_621));
INVX1 g42532(.A (n_621), .Y (n_838));
INVX1 g42249(.A (u10_mem_b1_b_120 ), .Y (n_6526));
INVX1 g42539(.A (u11_mem_b2_b ), .Y (n_419));
INVX1 g43110(.A (u11_mem_b3_b_86 ), .Y (n_5508));
INVX1 g41912(.A (u5_wp_b1_b ), .Y (n_734));
NAND2X1 g45819(.A (n_12537), .B (n_12538), .Y (n_12539));
OAI21X1 g45818(.A0 (n_5723), .A1 (n_7077), .B0 (n_6195), .Y(n_12533));
INVX1 g43114(.A (n_145), .Y (n_6134));
INVX1 g43117(.A (n_6824), .Y (n_6131));
AOI22X1 g40411(.A0 (u13_intm_r_b27_b ), .A1 (u13_ints_r_b27_b ), .B0(u13_intm_r_b28_b ), .B1 (u13_ints_r_b28_b ), .Y (n_731));
NAND2X1 g45812(.A (n_12389), .B (u4_mem_b0_b_94 ), .Y (n_12526));
NAND2X1 g39899(.A (u3_mem_b2_b ), .B (n_12619), .Y (n_2893));
OAI21X1 g45817(.A0 (n_12533), .A1 (n_12539), .B0 (n_10481), .Y(n_12543));
INVX1 g41910(.A (n_734), .Y (n_657));
NAND2X1 g45815(.A (n_3546), .B (u4_mem_b3_b_125 ), .Y (n_12529));
NAND2X1 g45814(.A (n_12087), .B (u4_mem_b2_b_32 ), .Y (n_12528));
NAND2X1 g39078(.A (u6_mem_b2_b_56 ), .B (n_3423), .Y (n_3468));
MX2X1 g34151(.A (u8_mem_b0_b_118 ), .B (n_3686), .S0 (n_7490), .Y(n_9378));
AOI21X1 g35598(.A0 (n_5932), .A1 (n_6121), .B0 (n_12604), .Y(n_7264));
AOI21X1 g35595(.A0 (n_5933), .A1 (n_5768), .B0 (n_7267), .Y (n_7127));
AOI21X1 g35594(.A0 (n_5934), .A1 (n_5769), .B0 (n_7267), .Y (n_7128));
AOI21X1 g35597(.A0 (n_6314), .A1 (n_6092), .B0 (n_7267), .Y (n_7265));
AOI21X1 g35596(.A0 (n_6819), .A1 (n_6130), .B0 (n_12145), .Y(n_7318));
AOI21X1 g35591(.A0 (n_6315), .A1 (n_5773), .B0 (n_7267), .Y (n_7266));
AOI21X1 g35590(.A0 (n_5937), .A1 (n_5774), .B0 (n_7267), .Y (n_7132));
AOI21X1 g35593(.A0 (n_5935), .A1 (n_5770), .B0 (n_12604), .Y(n_7129));
AOI21X1 g35592(.A0 (n_5936), .A1 (n_5771), .B0 (n_12604), .Y(n_7130));
INVX1 g36868(.A (n_6237), .Y (n_5722));
NAND4X1 g36869(.A (n_11646), .B (n_11647), .C (n_3166), .D (n_3532),.Y (n_6237));
AOI22X1 g40412(.A0 (u13_intm_r_b17_b ), .A1 (u13_ints_r_b17_b ), .B0(u13_intm_r_b18_b ), .B1 (u13_ints_r_b18_b ), .Y (n_576));
NAND2X1 g36860(.A (n_3925), .B (n_1248), .Y (n_5390));
NAND2X1 g36861(.A (n_1687), .B (n_3923), .Y (n_5389));
NAND2X1 g36862(.A (n_1572), .B (n_1571), .Y (n_4038));
NAND2X1 g36863(.A (n_3922), .B (n_1247), .Y (n_5388));
NAND2X1 g36864(.A (n_3921), .B (n_1245), .Y (n_5387));
INVX1 g36865(.A (n_6157), .Y (n_5723));
NAND4X1 g36866(.A (n_12004), .B (n_12005), .C (n_3336), .D (n_2450),.Y (n_6157));
NAND2X1 g36867(.A (n_2559), .B (n_3919), .Y (n_5386));
INVX1 g41918(.A (oc3_cfg_996), .Y (n_471));
INVX1 g41919(.A (u10_mem_b3_b_62 ), .Y (n_6565));
AOI22X1 g40413(.A0 (u13_intm_r_b21_b ), .A1 (u13_ints_r_b21_b ), .B0(u13_intm_r_b22_b ), .B1 (u13_ints_r_b22_b ), .Y (n_730));
NOR2X1 g39994(.A (n_2135), .B (n_2732), .Y (n_2211));
NAND2X1 g39844(.A (n_2344), .B (in_slt_422), .Y (n_2240));
NOR2X1 g40828(.A (n_6316), .B (u3_rp_b3_b ), .Y (n_664));
NOR2X1 g39997(.A (n_2218), .B (n_2712), .Y (n_1673));
NAND2X1 g39329(.A (u5_mem_b1_b ), .B (n_3236), .Y (n_11495));
OR2X1 g35319(.A (n_11563), .B (in_valid_s_b0_b ), .Y (n_7480));
NOR2X1 g39996(.A (n_2477), .B (n_2686), .Y (n_2209));
INVX1 g39322(.A (n_4769), .Y (n_3275));
NAND2X1 g39323(.A (in_slt_413), .B (n_2368), .Y (n_4769));
NAND2X1 g39320(.A (u7_mem_b2_b_30 ), .B (n_12654), .Y (n_3277));
AOI21X1 g38178(.A0 (u4_mem_b2_b_34 ), .A1 (n_4439), .B0 (n_2372), .Y(n_4410));
OAI21X1 g33568(.A0 (n_4409), .A1 (n_8333), .B0 (n_7989), .Y (n_8268));
NAND2X1 g34249(.A (u8_mem_b3_b_141 ), .B (n_7976), .Y (n_8153));
MX2X1 g38609(.A (u4_mem_b0_b_102 ), .B (wb_din_672), .S0 (n_3765), .Y(n_3799));
AOI21X1 g38179(.A0 (u4_mem_b2_b_35 ), .A1 (n_4439), .B0 (n_2095), .Y(n_4409));
NAND2X1 g34242(.A (u8_mem_b3_b_134 ), .B (n_7976), .Y (n_8163));
NAND2X1 g34243(.A (u8_mem_b3_b_135 ), .B (n_7976), .Y (n_8162));
OAI21X1 g33560(.A0 (n_4419), .A1 (n_8333), .B0 (n_7997), .Y (n_8277));
NAND2X1 g34241(.A (u3_mem_b1_b_62 ), .B (n_8101), .Y (n_8164));
NAND2X1 g34246(.A (u8_mem_b3_b_138 ), .B (n_7976), .Y (n_8157));
NAND2X1 g34247(.A (u8_mem_b3_b_139 ), .B (n_7976), .Y (n_8156));
OAI21X1 g33564(.A0 (n_4414), .A1 (n_9336), .B0 (n_7993), .Y (n_8272));
NAND2X1 g34245(.A (u3_mem_b1_b_64 ), .B (n_8101), .Y (n_8158));
NAND2X1 g39324(.A (u6_mem_b1_b_66 ), .B (n_4253), .Y (n_11716));
NAND3X1 g39325(.A (u5_mem_b0_b_92 ), .B (n_886), .C (n_1033), .Y(n_1319));
NOR2X1 g37531(.A (n_5313), .B (n_6649), .Y (n_4651));
OAI21X1 g37530(.A0 (n_1894), .A1 (u4_rp_b3_b ), .B0 (n_5466), .Y(n_5467));
NAND2X1 g37533(.A (n_5656), .B (n_4161), .Y (n_5244));
NOR2X1 g37532(.A (n_5304), .B (n_6649), .Y (n_4650));
NOR2X1 g37535(.A (n_5280), .B (n_6649), .Y (n_4649));
NAND2X1 g37534(.A (n_5656), .B (n_4193), .Y (n_5243));
NAND2X1 g37537(.A (n_5645), .B (n_3061), .Y (n_4648));
NOR2X1 g37536(.A (n_4767), .B (n_5371), .Y (n_3953));
NAND2X1 g37539(.A (n_635), .B (in_slt_742), .Y (n_1021));
NAND2X1 g37538(.A (n_5480), .B (n_2989), .Y (n_4647));
OAI21X1 g33621(.A0 (n_5027), .A1 (n_9290), .B0 (n_7921), .Y (n_9294));
OAI21X1 g33620(.A0 (n_5028), .A1 (n_9288), .B0 (n_7922), .Y (n_9296));
OAI21X1 g33623(.A0 (n_5025), .A1 (n_9288), .B0 (n_7919), .Y (n_9292));
OAI21X1 g33622(.A0 (n_5026), .A1 (n_9264), .B0 (n_7920), .Y (n_9293));
OAI21X1 g33625(.A0 (n_5022), .A1 (n_9288), .B0 (n_7917), .Y (n_9289));
OAI21X1 g33624(.A0 (n_5024), .A1 (n_9290), .B0 (n_7918), .Y (n_9291));
OAI21X1 g33627(.A0 (n_5018), .A1 (n_9235), .B0 (n_7915), .Y (n_9285));
OAI21X1 g33626(.A0 (n_5021), .A1 (n_9286), .B0 (n_7916), .Y (n_9287));
OAI21X1 g33629(.A0 (n_5016), .A1 (n_9202), .B0 (n_7913), .Y (n_9282));
OAI21X1 g33628(.A0 (n_5017), .A1 (n_9307), .B0 (n_7914), .Y (n_9283));
AOI22X1 g40418(.A0 (u13_intm_r_b11_b ), .A1 (u13_ints_r_b11_b ), .B0(u13_intm_r_b12_b ), .B1 (u13_ints_r_b12_b ), .Y (n_725));
NOR2X1 g39993(.A (n_2832), .B (n_2829), .Y (n_2830));
AOI21X1 g38175(.A0 (u4_mem_b2_b_32 ), .A1 (n_4439), .B0 (n_2066), .Y(n_4413));
AND2X1 g40901(.A (u10_rp_b1_b ), .B (n_403), .Y (n_2553));
AOI22X1 g40419(.A0 (u13_intm_r_b25_b ), .A1 (u13_ints_r_b25_b ), .B0(u13_intm_r_b26_b ), .B1 (u13_ints_r_b26_b ), .Y (n_577));
AOI21X1 g38529(.A0 (u4_mem_b1_b_65 ), .A1 (n_2470), .B0 (n_2481), .Y(n_4297));
AOI21X1 g38528(.A0 (u7_mem_b3_b ), .A1 (n_4961), .B0 (n_2890), .Y(n_4875));
AOI21X1 g38527(.A0 (u8_mem_b2_b_50 ), .A1 (n_4491), .B0 (n_1931), .Y(n_4298));
XOR2X1 g38526(.A (n_1443), .B (n_4961), .Y (n_4299));
AOI21X1 g38525(.A0 (u7_mem_b3_b_149 ), .A1 (n_4961), .B0 (n_3172), .Y(n_4876));
AOI21X1 g38524(.A0 (u7_mem_b3_b_130 ), .A1 (n_4961), .B0 (n_3446), .Y(n_4877));
AOI21X1 g38523(.A0 (u7_mem_b3_b_124 ), .A1 (n_5145), .B0 (n_3444), .Y(n_4878));
AOI21X1 g38522(.A0 (u7_mem_b3_b_151 ), .A1 (n_4961), .B0 (n_3015), .Y(n_4879));
AOI21X1 g38520(.A0 (u5_mem_b2_b_30 ), .A1 (n_4378), .B0 (n_2177), .Y(n_4300));
MX2X1 g33199(.A (u13_intm_r_b18_b ), .B (wb_din_678), .S0 (n_8519), .Y(n_8511));
MX2X1 g33198(.A (u13_intm_r_b17_b ), .B (wb_din_677), .S0 (n_8519), .Y(n_8512));
MX2X1 g33193(.A (u13_intm_r_b12_b ), .B (wb_din_672), .S0 (n_8519), .Y(n_8517));
MX2X1 g33192(.A (u13_intm_r_b11_b ), .B (wb_din_671), .S0 (n_8519), .Y(n_8518));
MX2X1 g33191(.A (u13_intm_r_b10_b ), .B (wb_din_670), .S0 (n_8519), .Y(n_8520));
MX2X1 g33190(.A (u13_intm_r_b0_b ), .B (wb_din), .S0 (n_8519), .Y(n_8521));
MX2X1 g33197(.A (u13_intm_r_b16_b ), .B (wb_din_676), .S0 (n_8519), .Y(n_8513));
MX2X1 g33196(.A (u13_intm_r_b15_b ), .B (wb_din_675), .S0 (n_8519), .Y(n_8514));
MX2X1 g33195(.A (u13_intm_r_b14_b ), .B (wb_din_674), .S0 (n_8519), .Y(n_8515));
MX2X1 g33194(.A (u13_intm_r_b13_b ), .B (wb_din_673), .S0 (n_8519), .Y(n_8516));
NAND2X1 g37129(.A (n_2498), .B (n_1706), .Y (n_3997));
AOI21X1 g38358(.A0 (u5_mem_b3_b_148 ), .A1 (n_5000), .B0 (n_3346), .Y(n_4979));
INVX1 g42788(.A (n_8567), .Y (n_942));
AOI21X1 g38359(.A0 (u5_mem_b3_b_149 ), .A1 (n_5000), .B0 (n_3123), .Y(n_4978));
INVX1 g42322(.A (u11_mem_b2_b_88 ), .Y (n_6454));
MX2X1 g38606(.A (u4_mem_b0_b ), .B (wb_din), .S0 (n_3765), .Y(n_3803));
AOI22X1 g37656(.A0 (u9_din_tmp_53), .A1 (n_2368), .B0 (in_slt_408),.B1 (n_3935), .Y (n_3938));
AOI22X1 g37657(.A0 (u9_din_tmp_54), .A1 (n_2368), .B0 (in_slt_409),.B1 (n_3935), .Y (n_3937));
INVX4 g41052(.A (n_1412), .Y (n_3236));
MX2X1 g38602(.A (u3_mem_b0_b_100 ), .B (wb_din_670), .S0 (n_3807), .Y(n_3809));
AOI22X1 g37651(.A0 (n_2502), .A1 (n_6847), .B0 (n_6928), .B1(n_1835), .Y (n_1709));
MX2X1 g38600(.A (u3_mem_b0_b_102 ), .B (wb_din_672), .S0 (n_3807), .Y(n_3812));
OAI21X1 g36668(.A0 (n_4587), .A1 (n_5183), .B0 (n_5772), .Y (n_5764));
AND2X1 g36669(.A (n_3967), .B (n_4685), .Y (n_5584));
OAI21X1 g36666(.A0 (n_5215), .A1 (n_5458), .B0 (n_6118), .Y (n_6119));
NAND2X1 g36667(.A (n_5557), .B (n_6091), .Y (n_6117));
NAND2X1 g36664(.A (n_5254), .B (n_3978), .Y (n_5765));
NAND2X1 g36665(.A (n_5538), .B (n_6091), .Y (n_6121));
OAI21X1 g36662(.A0 (n_4590), .A1 (n_4589), .B0 (n_5772), .Y (n_5768));
OAI21X1 g36663(.A0 (n_5167), .A1 (n_5166), .B0 (n_634), .Y (n_5767));
OAI21X1 g36660(.A0 (n_4581), .A1 (n_4591), .B0 (n_5772), .Y (n_5769));
OAI21X1 g36661(.A0 (n_5214), .A1 (n_5460), .B0 (n_6118), .Y (n_6122));
NOR2X1 g40136(.A (n_2790), .B (n_933), .Y (n_2098));
NAND2X1 g39656(.A (u7_mem_b2_b_29 ), .B (n_12645), .Y (n_3029));
NOR2X1 g30711(.A (n_10822), .B (n_5839), .Y (n_11008));
NOR2X1 g30712(.A (n_10775), .B (n_11136), .Y (n_10960));
NOR2X1 g30713(.A (n_10661), .B (n_11136), .Y (n_10959));
AND2X1 g30714(.A (n_10140), .B (n_2343), .Y (n_10807));
AND2X1 g30715(.A (n_10139), .B (n_9833), .Y (n_10806));
OAI21X1 g30716(.A0 (n_5840), .A1 (n_9615), .B0 (n_9614), .Y (n_9616));
OAI21X1 g30717(.A0 (n_5832), .A1 (n_9660), .B0 (n_9659), .Y (n_9661));
OAI21X1 g30718(.A0 (n_5438), .A1 (n_9612), .B0 (n_9611), .Y (n_9613));
OAI21X1 g30719(.A0 (n_5828), .A1 (n_9657), .B0 (n_9656), .Y (n_9658));
NAND2X1 g41059(.A (n_4683), .B (n_667), .Y (n_1153));
OR2X1 g41749(.A (n_523), .B (n_11612), .Y (n_829));
INVX1 g42200(.A (ic1_cfg_1036), .Y (n_625));
NAND2X1 g39657(.A (n_2344), .B (in_slt_432), .Y (n_2270));
NAND2X1 g41453(.A (u8_wp_b0_b ), .B (u8_wp_b1_b ), .Y (n_507));
INVX2 g41452(.A (n_507), .Y (n_982));
INVX4 g41450(.A (n_982), .Y (n_3879));
MX2X1 g36008(.A (n_6547), .B (n_6625), .S0 (n_6649), .Y (n_6626));
MX2X1 g36009(.A (n_6925), .B (n_6924), .S0 (n_5371), .Y (n_6926));
MX2X1 g36002(.A (n_6633), .B (n_6576), .S0 (n_5341), .Y (n_6634));
MX2X1 g36003(.A (n_6933), .B (n_6916), .S0 (n_930), .Y (n_6934));
MX2X1 g36000(.A (n_6635), .B (n_6582), .S0 (n_6898), .Y (n_6636));
MX2X1 g36001(.A (n_6935), .B (n_6952), .S0 (n_6898), .Y (n_6936));
MX2X1 g36006(.A (n_6928), .B (n_6927), .S0 (n_6898), .Y (n_6929));
MX2X1 g36007(.A (n_6628), .B (n_6560), .S0 (n_6898), .Y (n_6629));
MX2X1 g36004(.A (n_6630), .B (n_6573), .S0 (n_5341), .Y (n_6631));
MX2X1 g36005(.A (n_6931), .B (n_6896), .S0 (n_930), .Y (n_6932));
NOR2X1 g39654(.A (n_4996), .B (n_2765), .Y (n_3031));
NAND2X1 g45664(.A (n_11846), .B (n_11843), .Y (n_12354));
NOR2X1 g39998(.A (n_2827), .B (n_2864), .Y (n_2828));
NAND2X1 g39655(.A (n_11804), .B (u8_mem_b0_b_110 ), .Y (n_3030));
INVX1 g42327(.A (n_1921), .Y (n_1184));
INVX2 g41753(.A (n_835), .Y (n_1103));
NOR2X1 g39652(.A (n_5059), .B (n_2772), .Y (n_3035));
NAND2X1 g34747(.A (u7_mem_b1_b_66 ), .B (n_7651), .Y (n_7687));
NAND2X1 g34746(.A (u7_mem_b1_b_65 ), .B (n_7651), .Y (n_7688));
NAND2X1 g34745(.A (u7_mem_b1_b_64 ), .B (n_7651), .Y (n_7689));
NAND2X1 g34744(.A (u7_mem_b1_b_63 ), .B (n_7651), .Y (n_7690));
NAND2X1 g34743(.A (u7_mem_b1_b_62 ), .B (n_7651), .Y (n_7691));
NAND2X1 g34742(.A (u7_mem_b1_b_89 ), .B (n_7651), .Y (n_7692));
NAND2X1 g34741(.A (u7_mem_b1_b_61 ), .B (n_7651), .Y (n_7693));
NAND2X1 g34740(.A (u3_mem_b1_b_83 ), .B (n_8101), .Y (n_7694));
NAND2X1 g34749(.A (u7_mem_b1_b_68 ), .B (n_7651), .Y (n_7685));
OR2X1 g35292(.A (n_324), .B (n_11827), .Y (n_9579));
NAND2X1 g35293(.A (out_slt_24), .B (n_11827), .Y (n_9470));
OR2X1 g35290(.A (n_36), .B (n_11827), .Y (n_9472));
NAND2X1 g35291(.A (out_slt_25), .B (n_11827), .Y (n_9471));
OAI21X1 g35920(.A0 (n_5545), .A1 (n_7080), .B0 (n_5817), .Y (n_6987));
OR2X1 g35297(.A (n_5839), .B (n_11827), .Y (n_8671));
INVX1 g35294(.A (n_11841), .Y (n_9480));
OAI21X1 g35923(.A0 (n_6084), .A1 (n_11934), .B0 (n_6181), .Y(n_7177));
NAND2X1 g39249(.A (u4_mem_b1_b_62 ), .B (n_12259), .Y (n_4208));
NOR2X1 g39248(.A (u9_mem_b2_b_106 ), .B (n_1221), .Y (n_1222));
INVX1 g35298(.A (n_8670), .Y (n_9479));
INVX1 g35299(.A (n_7542), .Y (n_8670));
OAI21X1 g35928(.A0 (n_5675), .A1 (n_7063), .B0 (n_5816), .Y (n_7069));
OR2X1 g39651(.A (n_7256), .B (n_6821), .Y (n_2271));
NAND2X1 g34523(.A (u5_mem_b2_b ), .B (n_7870), .Y (n_7904));
NAND2X1 g34522(.A (u7_mem_b1_b_90 ), .B (n_7651), .Y (n_7906));
NAND2X1 g34521(.A (u5_mem_b1_b_68 ), .B (n_7870), .Y (n_7907));
NAND2X1 g34520(.A (u5_mem_b1_b_67 ), .B (n_7870), .Y (n_7908));
NAND2X1 g34527(.A (u5_mem_b2_b_41 ), .B (n_7870), .Y (n_7900));
NAND2X1 g34526(.A (u5_mem_b2_b_40 ), .B (n_7870), .Y (n_7901));
NAND2X1 g34525(.A (u5_mem_b2_b_39 ), .B (n_7870), .Y (n_7902));
NAND2X1 g34524(.A (u5_mem_b2_b_38 ), .B (n_7870), .Y (n_7903));
MX2X1 g31281(.A (n_6387), .B (n_6386), .S0 (n_10137), .Y (n_10136));
NAND2X1 g34529(.A (u5_mem_b2_b_43 ), .B (n_7870), .Y (n_7898));
NAND2X1 g34528(.A (u5_mem_b2_b_42 ), .B (n_7870), .Y (n_7899));
MX2X1 g38604(.A (u7_mem_b0_b_101 ), .B (wb_din_671), .S0 (n_913), .Y(n_3806));
INVX2 g41722(.A (n_813), .Y (n_1106));
NOR2X1 g29980(.A (n_10406), .B (dma_ack_i_b5_b), .Y (n_11122));
AOI21X1 g35436(.A0 (n_1560), .A1 (n_2302), .B0 (n_3941), .Y (n_5447));
AOI21X1 g35437(.A0 (n_1234), .A1 (n_2513), .B0 (n_2569), .Y (n_4848));
AOI21X1 g35434(.A0 (n_6959), .A1 (n_4741), .B0 (n_7353), .Y (n_7339));
AOI21X1 g35435(.A0 (n_1558), .A1 (n_2368), .B0 (n_2570), .Y (n_4850));
AOI21X1 g35432(.A0 (n_6962), .A1 (n_4697), .B0 (n_7353), .Y (n_7341));
AOI21X1 g35433(.A0 (n_6961), .A1 (n_4695), .B0 (n_7353), .Y (n_7340));
AOI21X1 g35430(.A0 (n_6964), .A1 (n_4702), .B0 (n_7353), .Y (n_7343));
AOI21X1 g35431(.A0 (n_6963), .A1 (n_4698), .B0 (n_7353), .Y (n_7342));
NOR2X1 g35438(.A (n_7025), .B (n_1133), .Y (n_7028));
NOR2X1 g35439(.A (n_7019), .B (n_7022), .Y (n_7027));
CLKBUFX1 g32807(.A (n_9633), .Y (n_9681));
INVX4 g32805(.A (n_9681), .Y (n_10738));
NOR2X1 g35810(.A (n_694), .B (n_6752), .Y (n_6740));
NAND2X1 g36480(.A (n_5867), .B (n_5876), .Y (n_5868));
NOR2X1 g40007(.A (n_2025), .B (n_2782), .Y (n_2203));
NOR2X1 g40005(.A (n_2477), .B (n_2782), .Y (n_2205));
NOR2X1 g40004(.A (n_2790), .B (n_1985), .Y (n_1826));
NOR2X1 g40001(.A (n_821), .B (n_2732), .Y (n_2208));
NOR2X1 g40000(.A (n_2736), .B (n_2782), .Y (n_2824));
NOR2X1 g40009(.A (n_1016), .B (n_2684), .Y (n_2822));
NOR2X1 g40008(.A (n_2827), .B (n_2763), .Y (n_2823));
OR2X1 g41729(.A (wb_addr_i_b31_b), .B (wb_addr_i_b29_b), .Y (n_421));
NOR2X1 g40002(.A (n_2470), .B (n_2716), .Y (n_2207));
NOR2X1 g41728(.A (u11_rp_b2_b ), .B (u11_wp_b3_b ), .Y (n_522));
INVX1 g42242(.A (u9_mem_b0_b_168 ), .Y (n_174));
NAND2X1 g39377(.A (u8_mem_b1_b_67 ), .B (n_12295), .Y (n_11448));
INVX1 g42813(.A (oc4_cfg_1009), .Y (n_454));
OR2X1 g41505(.A (n_11597), .B (n_1124), .Y (n_1126));
MX2X1 g37276(.A (u9_mem_b1_b_144 ), .B (n_4749), .S0 (n_5730), .Y(n_4750));
MX2X1 g37277(.A (u10_mem_b2_b_116 ), .B (n_5284), .S0 (n_5341), .Y(n_5342));
MX2X1 g37274(.A (u10_mem_b2_b_115 ), .B (n_4751), .S0 (n_5341), .Y(n_4752));
AOI21X1 g37275(.A0 (n_5488), .A1 (n_6649), .B0 (n_4654), .Y (n_5489));
AOI21X1 g37272(.A0 (n_5345), .A1 (n_5371), .B0 (n_3960), .Y (n_5346));
AOI21X1 g37273(.A0 (n_5343), .A1 (n_5371), .B0 (n_3950), .Y (n_5344));
AOI21X1 g37270(.A0 (n_5347), .A1 (n_5371), .B0 (n_3961), .Y (n_5348));
MX2X1 g37271(.A (u9_mem_b1_b_142 ), .B (n_4753), .S0 (n_4783), .Y(n_4754));
MX2X1 g37278(.A (u10_mem_b2_b_118 ), .B (n_5339), .S0 (n_5424), .Y(n_5340));
MX2X1 g37279(.A (u9_mem_b2_b_108 ), .B (n_4747), .S0 (n_6898), .Y(n_4748));
INVX2 g41202(.A (n_12172), .Y (n_1845));
INVX4 g41200(.A (n_1845), .Y (n_4253));
INVX1 g42247(.A (u11_mem_b3_b_75 ), .Y (n_5582));
BUFX3 g41600(.A (n_5102), .Y (n_5106));
INVX4 g40917(.A (n_1163), .Y (n_5312));
INVX1 g40916(.A (n_932), .Y (n_1163));
OAI21X1 g31058(.A0 (n_4766), .A1 (n_10679), .B0 (n_9980), .Y(n_10805));
OAI21X1 g31059(.A0 (n_4780), .A1 (n_10679), .B0 (n_9979), .Y(n_10667));
NAND2X1 g31728(.A (n_5524), .B (n_10391), .Y (n_10347));
NAND2X1 g31729(.A (n_5508), .B (n_10385), .Y (n_10346));
OAI21X1 g31054(.A0 (n_5291), .A1 (n_10679), .B0 (n_9984), .Y(n_10672));
OAI21X1 g31055(.A0 (n_5289), .A1 (n_10450), .B0 (n_9983), .Y(n_10671));
OAI21X1 g31056(.A0 (n_5288), .A1 (n_10450), .B0 (n_9982), .Y(n_10670));
OAI21X1 g31057(.A0 (n_5356), .A1 (n_10450), .B0 (n_9981), .Y(n_10669));
OAI21X1 g31050(.A0 (n_5297), .A1 (n_10820), .B0 (n_10360), .Y(n_10860));
NAND2X1 g31723(.A (n_5496), .B (n_10376), .Y (n_10352));
OAI21X1 g31052(.A0 (n_5301), .A1 (n_10820), .B0 (n_10359), .Y(n_10859));
OAI21X1 g31053(.A0 (n_4746), .A1 (n_10679), .B0 (n_9985), .Y(n_10673));
NAND2X1 g34379(.A (u4_mem_b1_b_63 ), .B (n_7984), .Y (n_8024));
NAND2X1 g34748(.A (u7_mem_b1_b_67 ), .B (n_7651), .Y (n_7686));
AOI21X1 g33388(.A0 (n_8660), .A1 (n_1146), .B0 (n_1007), .Y (n_9507));
AOI21X1 g33389(.A0 (n_1309), .A1 (n_7480), .B0 (n_1260), .Y (n_8484));
AOI21X1 g33386(.A0 (n_8664), .A1 (n_1356), .B0 (n_1023), .Y (n_9509));
AOI21X1 g33387(.A0 (n_8662), .A1 (n_1101), .B0 (n_1008), .Y (n_9508));
AOI21X1 g33384(.A0 (n_8669), .A1 (n_1302), .B0 (n_1010), .Y (n_9511));
AOI21X1 g33385(.A0 (n_8666), .A1 (n_1373), .B0 (n_1009), .Y (n_9510));
NOR2X1 g33382(.A (n_5631), .B (u2_bit_clk_e), .Y (n_6065));
AOI21X1 g33383(.A0 (n_8671), .A1 (n_1375), .B0 (n_1021), .Y (n_9512));
INVX1 g33380(.A (n_9513), .Y (n_9564));
NOR2X1 g33381(.A (n_7536), .B (u14_u7_en_out_l2), .Y (n_9513));
INVX4 g40515(.A (wb_din_671), .Y (n_2716));
NAND2X1 g34373(.A (u4_mem_b1_b_88 ), .B (n_7984), .Y (n_8029));
OAI21X1 g33410(.A0 (n_3851), .A1 (n_8464), .B0 (n_7838), .Y (n_8465));
NAND2X1 g34371(.A (u4_mem_b1_b_86 ), .B (n_7984), .Y (n_8031));
AOI21X1 g35618(.A0 (n_5830), .A1 (n_6820), .B0 (n_7256), .Y (n_7311));
OAI21X1 g33416(.A0 (n_3884), .A1 (n_8433), .B0 (n_8160), .Y (n_8456));
AOI21X1 g30887(.A0 (n_11621), .A1 (n_11622), .B0 (n_11030), .Y(n_11031));
NAND2X1 g39552(.A (n_2491), .B (u7_mem_b0_b_97 ), .Y (n_1809));
OAI21X1 g33417(.A0 (n_5153), .A1 (n_8911), .B0 (n_7618), .Y (n_8455));
AOI21X1 g35616(.A0 (n_5919), .A1 (n_6106), .B0 (n_12640), .Y(n_7247));
NAND2X1 g34374(.A (u4_mem_b1_b_61 ), .B (n_7984), .Y (n_8028));
AOI21X1 g30889(.A0 (n_11731), .A1 (n_11732), .B0 (n_11043), .Y(n_11028));
OAI21X1 g33415(.A0 (n_3845), .A1 (n_8457), .B0 (n_8162), .Y (n_8458));
NAND2X1 g36495(.A (n_12171), .B (n_6816), .Y (n_6789));
NAND2X1 g36494(.A (n_12531), .B (n_6790), .Y (n_6791));
NAND2X1 g36497(.A (n_6233), .B (n_6773), .Y (n_6234));
AOI21X1 g35615(.A0 (n_5920), .A1 (n_6223), .B0 (n_7256), .Y (n_7248));
NAND2X1 g36491(.A (n_6816), .B (n_5855), .Y (n_5856));
NAND2X1 g36490(.A (n_6237), .B (n_12531), .Y (n_6238));
NAND2X1 g36492(.A (n_6235), .B (n_12115), .Y (n_6236));
INVX4 g40652(.A (wb_din_687), .Y (n_2763));
NAND2X1 g36499(.A (n_6816), .B (n_5851), .Y (n_5852));
NAND2X1 g36498(.A (n_6786), .B (n_6816), .Y (n_6787));
INVX1 g43023(.A (u11_mem_b1_b_128 ), .Y (n_6519));
NAND2X1 g39589(.A (u8_mem_b1_b_78 ), .B (n_12291), .Y (n_3078));
AOI21X1 g35609(.A0 (n_6826), .A1 (n_6111), .B0 (n_7256), .Y (n_7315));
AOI21X1 g35608(.A0 (n_6823), .A1 (n_6112), .B0 (n_7256), .Y (n_7316));
AOI21X1 g30899(.A0 (n_11637), .A1 (n_11638), .B0 (n_11025), .Y(n_11019));
AOI21X1 g30898(.A0 (n_11992), .A1 (n_11993), .B0 (n_11036), .Y(n_11020));
AOI21X1 g35605(.A0 (n_5926), .A1 (n_6116), .B0 (n_7256), .Y (n_7257));
NOR2X1 g30896(.A (n_10973), .B (n_11128), .Y (n_11129));
NOR2X1 g30895(.A (n_10974), .B (n_11128), .Y (n_11130));
AOI21X1 g30894(.A0 (n_12016), .A1 (n_12017), .B0 (n_5839), .Y(n_11022));
AOI21X1 g30893(.A0 (n_11629), .A1 (n_11630), .B0 (n_11033), .Y(n_11023));
AOI21X1 g30892(.A0 (n_11735), .A1 (n_11736), .B0 (n_5839), .Y(n_11024));
AOI21X1 g30891(.A0 (n_11625), .A1 (n_11626), .B0 (n_11025), .Y(n_11026));
AOI21X1 g30890(.A0 (n_11733), .A1 (n_11734), .B0 (n_11043), .Y(n_11027));
AOI22X1 g37834(.A0 (n_2344), .A1 (in_slt_436), .B0 (n_2302), .B1(in_slt_424), .Y (n_5418));
NAND2X1 g37835(.A (n_3016), .B (n_3360), .Y (n_4580));
AOI22X1 g37344(.A0 (n_5277), .A1 (crac_out_876), .B0 (n_6972), .B1(oc3_cfg_1000), .Y (n_5268));
NAND2X1 g38825(.A (u4_mem_b3_b_146 ), .B (n_3556), .Y (n_3550));
INVX1 g42517(.A (n_469), .Y (n_4688));
INVX1 g42515(.A (oc0_cfg_969), .Y (n_498));
INVX1 g42248(.A (u10_mem_b2_b_114 ), .Y (n_2627));
INVX2 g42512(.A (u4_rp_b1_b ), .Y (n_551));
INVX1 g42511(.A (n_551), .Y (n_521));
NAND2X1 g38823(.A (u4_mem_b3_b_142 ), .B (n_3556), .Y (n_3551));
NOR2X1 g39726(.A (u10_mem_b1_b_132 ), .B (n_2364), .Y (n_2257));
NAND2X1 g39724(.A (u5_mem_b2_b_50 ), .B (n_12823), .Y (n_2250));
NAND2X1 g39725(.A (n_12204), .B (u6_mem_b0_b_121 ), .Y (n_2995));
INVX1 g39722(.A (n_5321), .Y (n_4138));
NAND2X1 g38820(.A (u4_mem_b3_b_124 ), .B (n_4258), .Y (n_4256));
NAND2X1 g39720(.A (n_11798), .B (u8_mem_b0_b_118 ), .Y (n_2997));
NAND2X1 g39721(.A (u3_mem_b2_b_44 ), .B (n_12619), .Y (n_2996));
NAND2X1 g38821(.A (u4_mem_b3_b_126 ), .B (n_3546), .Y (n_2634));
NAND2X1 g39058(.A (u3_mem_b1_b_68 ), .B (n_3316), .Y (n_12004));
INVX1 g39728(.A (n_4745), .Y (n_2994));
NAND2X1 g39729(.A (n_2302), .B (in_slt_427), .Y (n_4745));
NAND2X1 g36802(.A (n_1705), .B (n_1730), .Y (n_4050));
NAND2X1 g36803(.A (n_1729), .B (n_1726), .Y (n_4049));
NAND2X1 g36800(.A (n_1563), .B (n_1735), .Y (n_4052));
NAND2X1 g36801(.A (n_1734), .B (n_1699), .Y (n_4051));
NAND2X1 g36806(.A (n_1719), .B (n_1718), .Y (n_4046));
NAND2X1 g36807(.A (n_2508), .B (n_1858), .Y (n_4045));
NAND2X1 g36804(.A (n_1725), .B (n_1722), .Y (n_4048));
NAND2X1 g36805(.A (n_2501), .B (n_1720), .Y (n_4047));
AOI21X1 g38497(.A0 (u7_mem_b2_b_45 ), .A1 (n_4540), .B0 (n_2117), .Y(n_4314));
NAND2X1 g36808(.A (n_1717), .B (n_2505), .Y (n_4044));
NAND2X1 g36809(.A (n_1714), .B (n_1712), .Y (n_4043));
AOI21X1 g38496(.A0 (u7_mem_b2_b_43 ), .A1 (n_4509), .B0 (n_2185), .Y(n_4315));
NAND2X1 g39243(.A (n_4560), .B (in_slt_457), .Y (n_5298));
INVX1 g39242(.A (n_5298), .Y (n_4209));
NAND2X1 g38828(.A (u3_mem_b3_b_130 ), .B (n_2463), .Y (n_2450));
NOR2X1 g39245(.A (n_3332), .B (n_2720), .Y (n_3344));
NOR2X1 g36522(.A (o4_status), .B (n_5831), .Y (n_5832));
INVX8 g41609(.A (n_1475), .Y (n_3486));
NOR2X1 g39244(.A (u10_mem_b1_b_136 ), .B (n_2364), .Y (n_2341));
OAI21X1 g35922(.A0 (n_5685), .A1 (n_7077), .B0 (n_6193), .Y (n_7076));
NOR2X1 g41403(.A (u9_rp_b2_b ), .B (u9_wp_b3_b ), .Y (n_478));
NAND2X1 g39246(.A (u5_mem_b2_b_30 ), .B (n_12823), .Y (n_11443));
INVX4 g41550(.A (n_12621), .Y (n_2419));
INVX1 g42509(.A (n_761), .Y (n_1923));
NOR2X1 g41556(.A (n_693), .B (n_942), .Y (n_741));
AND2X1 g41557(.A (n_699), .B (n_872), .Y (n_7531));
INVX1 g41999(.A (u9_mem_b1_b_136 ), .Y (n_204));
INVX1 g41992(.A (n_667), .Y (n_4706));
INVX1 g41993(.A (ic2_cfg_1046), .Y (n_667));
INVX1 g41990(.A (u11_mem_b0_b_180 ), .Y (n_1581));
INVX1 g41991(.A (u11_mem_b0_b_162 ), .Y (n_6366));
INVX1 g41996(.A (u10_mem_b2_b_112 ), .Y (n_2549));
INVX1 g42974(.A (u9_mem_b2_b_109 ), .Y (n_198));
NOR2X1 g45651(.A (n_1374), .B (n_11507), .Y (n_12334));
INVX1 g41873(.A (u9_mem_b0_b_171 ), .Y (n_1738));
OAI21X1 g33544(.A0 (n_4436), .A1 (n_8333), .B0 (n_8013), .Y (n_8296));
OAI21X1 g33545(.A0 (n_4435), .A1 (n_8318), .B0 (n_8012), .Y (n_8295));
OAI21X1 g33814(.A0 (n_4901), .A1 (n_9055), .B0 (n_7713), .Y (n_9056));
OAI21X1 g33547(.A0 (n_4432), .A1 (n_8333), .B0 (n_8010), .Y (n_8293));
NAND2X1 g34260(.A (u3_mem_b2_b_39 ), .B (n_8141), .Y (n_8142));
OAI21X1 g33541(.A0 (n_4440), .A1 (n_8318), .B0 (n_8016), .Y (n_8300));
OAI21X1 g33810(.A0 (n_4904), .A1 (n_9055), .B0 (n_7718), .Y (n_9062));
OAI21X1 g33811(.A0 (n_4929), .A1 (n_9055), .B0 (n_7717), .Y (n_9061));
NAND2X1 g39370(.A (u5_mem_b2_b_54 ), .B (n_12823), .Y (n_2316));
INVX1 g45652(.A (n_12335), .Y (n_12336));
NAND2X1 g34268(.A (u3_mem_b2_b_42 ), .B (n_8141), .Y (n_8132));
NAND2X1 g34269(.A (u3_mem_b2_b_43 ), .B (n_8101), .Y (n_8131));
OAI21X1 g33818(.A0 (n_5083), .A1 (n_9034), .B0 (n_7707), .Y (n_9049));
OAI21X1 g33819(.A0 (n_4991), .A1 (n_8981), .B0 (n_7706), .Y (n_9048));
NAND2X1 g39906(.A (u5_mem_b1_b_80 ), .B (n_3239), .Y (n_2888));
NOR2X1 g40348(.A (n_2767), .B (n_2057), .Y (n_1946));
INVX1 g37049(.A (n_5541), .Y (n_5542));
MX2X1 g38728(.A (u7_mem_b0_b_120 ), .B (wb_din_690), .S0 (n_3622), .Y(n_3613));
AOI21X1 g38099(.A0 (u8_mem_b2_b_30 ), .A1 (n_4491), .B0 (n_2002), .Y(n_4479));
AOI21X1 g38016(.A0 (u3_mem_b2_b_39 ), .A1 (n_4533), .B0 (n_2075), .Y(n_4534));
INVX1 g37045(.A (n_6204), .Y (n_5687));
NAND4X1 g37044(.A (n_4247), .B (n_2200), .C (n_4196), .D (n_1395), .Y(n_6763));
NAND4X1 g37047(.A (n_4204), .B (n_2289), .C (n_2945), .D (n_1531), .Y(n_6228));
NAND4X1 g37046(.A (n_4210), .B (n_1499), .C (n_3277), .D (n_1275), .Y(n_6204));
NAND4X1 g37041(.A (n_4125), .B (n_2331), .C (n_2956), .D (n_1533), .Y(n_6207));
INVX1 g37043(.A (n_6763), .Y (n_6072));
NAND2X1 g37514(.A (n_5656), .B (n_4238), .Y (n_5245));
OAI21X1 g33609(.A0 (n_5042), .A1 (n_9286), .B0 (n_7936), .Y (n_9312));
OAI21X1 g33608(.A0 (n_5043), .A1 (n_9307), .B0 (n_7938), .Y (n_9313));
OAI21X1 g33603(.A0 (n_4384), .A1 (n_8856), .B0 (n_8132), .Y (n_9318));
OAI21X1 g33602(.A0 (n_5064), .A1 (n_9349), .B0 (n_7950), .Y (n_9319));
OAI21X1 g33601(.A0 (n_5065), .A1 (n_9349), .B0 (n_7951), .Y (n_9320));
OAI21X1 g33600(.A0 (n_5067), .A1 (n_9326), .B0 (n_7952), .Y (n_9321));
OAI21X1 g33607(.A0 (n_5023), .A1 (n_9307), .B0 (n_7939), .Y (n_9314));
OAI21X1 g33606(.A0 (n_5046), .A1 (n_9307), .B0 (n_7941), .Y (n_9315));
OAI21X1 g33605(.A0 (n_5047), .A1 (n_9286), .B0 (n_7942), .Y (n_9316));
OAI21X1 g33604(.A0 (n_5049), .A1 (n_9286), .B0 (n_7943), .Y (n_9317));
NAND2X1 g36877(.A (n_2551), .B (n_2548), .Y (n_4818));
NOR2X1 g39068(.A (n_2744), .B (n_1488), .Y (n_1502));
NAND2X1 g45760(.A (n_12479), .B (n_12482), .Y (n_12483));
NOR2X1 g37494(.A (n_4749), .B (n_5371), .Y (n_3963));
INVX1 g36872(.A (n_6244), .Y (n_5721));
AOI21X1 g38549(.A0 (u8_mem_b1_b_79 ), .A1 (n_4387), .B0 (n_1956), .Y(n_4283));
AOI21X1 g38548(.A0 (u8_mem_b1_b_78 ), .A1 (n_4387), .B0 (n_2122), .Y(n_4284));
NAND2X1 g36871(.A (n_1686), .B (n_1683), .Y (n_4037));
AOI21X1 g38541(.A0 (u8_mem_b1_b_88 ), .A1 (n_4502), .B0 (n_1987), .Y(n_4290));
AOI21X1 g38540(.A0 (u8_mem_b2_b_48 ), .A1 (n_4491), .B0 (n_2176), .Y(n_4291));
AOI21X1 g38543(.A0 (u8_mem_b3_b_133 ), .A1 (n_3879), .B0 (n_1556), .Y(n_3842));
AOI21X1 g38542(.A0 (u5_mem_b2_b_51 ), .A1 (n_4370), .B0 (n_1936), .Y(n_4289));
AOI21X1 g38545(.A0 (u8_mem_b1_b_72 ), .A1 (n_4387), .B0 (n_2119), .Y(n_4287));
AOI21X1 g38544(.A0 (u8_mem_b1_b_70 ), .A1 (n_4387), .B0 (n_1965), .Y(n_4288));
AOI21X1 g38547(.A0 (u8_mem_b1_b_76 ), .A1 (n_4502), .B0 (n_2202), .Y(n_4285));
AOI21X1 g38546(.A0 (u8_mem_b1_b_74 ), .A1 (n_4502), .B0 (n_1960), .Y(n_4286));
NAND2X1 g39061(.A (n_12825), .B (u3_mem_b0_b_114 ), .Y (n_3482));
NOR2X1 g40346(.A (n_2043), .B (n_2763), .Y (n_1948));
NAND2X1 g39060(.A (n_3252), .B (u7_mem_b0_b_110 ), .Y (n_3483));
NOR2X1 g40347(.A (n_2169), .B (n_2691), .Y (n_1947));
OAI21X1 g45779(.A0 (n_12499), .A1 (n_12500), .B0 (n_12504), .Y(n_12505));
NAND2X1 g32635(.A (n_370), .B (n_9947), .Y (n_12043));
NAND2X1 g32634(.A (n_380), .B (n_9947), .Y (n_11538));
NAND2X1 g32637(.A (n_391), .B (n_9943), .Y (n_11981));
NAND2X1 g32636(.A (n_351), .B (n_9947), .Y (n_11951));
AOI21X1 g32631(.A0 (n_6808), .A1 (n_6806), .B0 (n_10787), .Y(n_9941));
NAND2X1 g32630(.A (n_361), .B (n_9943), .Y (n_12013));
NAND2X1 g32633(.A (n_373), .B (n_9943), .Y (n_11536));
AOI21X1 g32632(.A0 (n_6804), .A1 (n_6801), .B0 (n_10787), .Y(n_9940));
NAND2X1 g32639(.A (u10_wp_b2_b ), .B (n_9564), .Y (n_9752));
NAND2X1 g32638(.A (n_394), .B (n_9947), .Y (n_12007));
NOR2X1 g39067(.A (n_2716), .B (n_1488), .Y (n_1435));
NAND2X1 g39066(.A (u8_mem_b2_b_35 ), .B (n_2362), .Y (n_2363));
NAND2X1 g36648(.A (n_5261), .B (n_2580), .Y (n_5782));
NAND2X1 g36649(.A (n_5260), .B (n_2579), .Y (n_5781));
NAND2X1 g36398(.A (n_5803), .B (n_2567), .Y (n_5906));
NAND2X1 g36399(.A (n_6250), .B (n_2567), .Y (n_6277));
OR2X1 g35462(.A (n_11762), .B (n_630), .Y (n_7441));
OAI21X1 g36640(.A0 (n_4606), .A1 (n_5218), .B0 (u4_rp_b0_b ), .Y(n_6124));
NAND2X1 g36393(.A (n_6184), .B (n_6316), .Y (n_6282));
NAND2X1 g36390(.A (n_5811), .B (n_2567), .Y (n_5909));
MX2X1 g31163(.A (n_6590), .B (n_6588), .S0 (n_9676), .Y (n_10228));
NAND2X1 g36396(.A (n_5809), .B (n_2567), .Y (n_5907));
NAND2X1 g36397(.A (n_11895), .B (n_6316), .Y (n_6278));
NAND2X1 g36394(.A (n_11898), .B (n_6316), .Y (n_6280));
NAND2X1 g36395(.A (n_6172), .B (n_6316), .Y (n_6279));
INVX1 g42369(.A (oc1_cfg_976), .Y (n_283));
NAND2X1 g38897(.A (u6_mem_b3_b_140 ), .B (n_2419), .Y (n_2417));
NAND2X1 g38896(.A (n_393), .B (n_831), .Y (n_3944));
NAND2X1 g38895(.A (u6_mem_b3_b_152 ), .B (n_2465), .Y (n_2418));
NAND2X1 g38894(.A (u6_mem_b3_b_138 ), .B (n_2419), .Y (n_2420));
NAND2X1 g38893(.A (u6_mem_b3_b_150 ), .B (n_2465), .Y (n_2421));
NAND2X1 g38891(.A (u6_mem_b3_b_136 ), .B (n_2419), .Y (n_2423));
NAND2X1 g38890(.A (u6_mem_b3_b_134 ), .B (n_2419), .Y (n_2424));
AOI22X1 g37820(.A0 (n_1756), .A1 (n_1615), .B0 (n_1614), .B1(n_1643), .Y (n_1616));
NAND2X1 g38898(.A (u6_mem_b3_b_122 ), .B (n_12622), .Y (n_2416));
MX2X1 g36024(.A (n_6906), .B (n_6905), .S0 (n_6908), .Y (n_6907));
MX2X1 g36025(.A (n_6018), .B (n_6017), .S0 (n_5341), .Y (n_6019));
MX2X1 g36027(.A (n_6599), .B (n_6598), .S0 (n_6594), .Y (n_6600));
MX2X1 g36020(.A (n_6916), .B (n_6915), .S0 (n_6908), .Y (n_6917));
MX2X1 g36021(.A (n_6021), .B (n_6003), .S0 (n_5341), .Y (n_6022));
MX2X1 g36022(.A (n_6913), .B (n_6912), .S0 (n_6908), .Y (n_6914));
MX2X1 g36023(.A (n_6927), .B (n_6909), .S0 (n_6908), .Y (n_6910));
INVX1 g41431(.A (n_3556), .Y (n_1894));
CLKBUFX3 g41430(.A (n_12743), .Y (n_3546));
NOR2X1 g39515(.A (n_3117), .B (n_2684), .Y (n_3129));
BUFX3 g41432(.A (n_12743), .Y (n_3556));
MX2X1 g36028(.A (n_6596), .B (n_6595), .S0 (n_6594), .Y (n_6597));
MX2X1 g36029(.A (n_6902), .B (n_6913), .S0 (n_6898), .Y (n_6903));
INVX1 g42304(.A (u7_wp_b1_b ), .Y (n_705));
INVX1 g42228(.A (u9_mem_b2_b_118 ), .Y (n_343));
AOI21X1 g38278(.A0 (u8_mem_b1_b_86 ), .A1 (n_4387), .B0 (n_2214), .Y(n_4382));
AOI22X1 g37773(.A0 (n_162), .A1 (n_1839), .B0 (n_5504), .B1 (n_1316),.Y (n_1663));
INVX1 g42305(.A (u9_mem_b3_b_85 ), .Y (n_5345));
CLKBUFX1 g45389(.A (n_11612), .Y (n_11597));
AOI21X1 g37772(.A0 (n_6424), .A1 (n_1831), .B0 (n_1211), .Y (n_1664));
AOI22X1 g37771(.A0 (n_1756), .A1 (n_6366), .B0 (n_6511), .B1(n_1643), .Y (n_1665));
NAND2X1 g37770(.A (n_3527), .B (n_2297), .Y (n_4587));
AOI22X1 g37777(.A0 (n_6415), .A1 (n_2530), .B0 (n_6633), .B1(n_2544), .Y (n_2532));
INVX8 g35160(.A (o8_we), .Y (n_7651));
AOI22X1 g37776(.A0 (n_6507), .A1 (n_1643), .B0 (n_6421), .B1(n_1831), .Y (n_1661));
AOI22X1 g37775(.A0 (u10_din_tmp_49), .A1 (n_2302), .B0 (n_3911), .B1(in_slt_428), .Y (n_2533));
XOR2X1 g40438(.A (n_1198), .B (n_2567), .Y (n_3992));
NOR2X1 g37135(.A (n_3560), .B (n_12823), .Y (n_5942));
NAND2X1 g34721(.A (u7_mem_b1_b_73 ), .B (n_7651), .Y (n_7716));
NAND2X1 g34720(.A (u7_mem_b1_b_72 ), .B (n_7651), .Y (n_7717));
NAND2X1 g34723(.A (u7_mem_b1_b_75 ), .B (n_7651), .Y (n_7713));
NAND2X1 g34722(.A (u7_mem_b1_b_74 ), .B (n_7651), .Y (n_7715));
NAND2X1 g34725(.A (u7_mem_b1_b_77 ), .B (n_7651), .Y (n_7710));
NOR2X1 g34896(.A (n_12838), .B (n_12837), .Y (n_7437));
NAND2X1 g34727(.A (u7_mem_b1_b_60 ), .B (n_7651), .Y (n_7707));
NAND2X1 g34726(.A (u7_mem_b1_b_78 ), .B (n_7651), .Y (n_7708));
NAND2X1 g34729(.A (u7_mem_b1_b_80 ), .B (n_7651), .Y (n_7705));
NAND2X1 g34728(.A (u7_mem_b1_b_79 ), .B (n_7651), .Y (n_7706));
NOR2X1 g34899(.A (n_7281), .B (n_3993), .Y (n_7435));
NOR2X1 g34898(.A (n_7282), .B (n_4796), .Y (n_7436));
INVX1 g42168(.A (u10_mem_b3_b_77 ), .Y (n_5363));
OAI21X1 g33066(.A0 (n_7122), .A1 (n_7065), .B0 (n_10483), .Y(n_11613));
NOR2X1 g39269(.A (n_3332), .B (n_2755), .Y (n_3333));
NAND2X1 g39268(.A (u8_mem_b2_b_31 ), .B (n_3334), .Y (n_12038));
NAND2X1 g39919(.A (n_11804), .B (u8_mem_b0_b_115 ), .Y (n_2876));
NOR2X1 g39918(.A (n_3486), .B (n_2782), .Y (n_2877));
NOR2X1 g39263(.A (n_5138), .B (n_2748), .Y (n_3338));
NAND2X1 g39262(.A (n_3339), .B (in_slt_437), .Y (n_5339));
INVX1 g39261(.A (n_5339), .Y (n_4206));
NAND2X1 g39260(.A (u8_mem_b2_b_44 ), .B (n_3334), .Y (n_12036));
NAND2X1 g39267(.A (u3_mem_b2_b_37 ), .B (n_12619), .Y (n_3336));
NAND2X1 g39266(.A (n_4560), .B (in_slt_449), .Y (n_5317));
INVX1 g39265(.A (n_5317), .Y (n_4205));
NOR2X1 g39264(.A (u10_mem_b1_b_119 ), .B (n_2364), .Y (n_2336));
MX2X1 g34099(.A (u7_mem_b0_b_113 ), .B (n_3569), .S0 (n_7493), .Y(n_8739));
MX2X1 g34098(.A (u7_mem_b0_b_112 ), .B (n_3641), .S0 (n_7493), .Y(n_9396));
MX2X1 g34093(.A (u7_mem_b0_b_108 ), .B (n_3564), .S0 (n_7493), .Y(n_8745));
MX2X1 g34092(.A (u7_mem_b0_b_107 ), .B (n_3644), .S0 (n_7493), .Y(n_8747));
MX2X1 g34091(.A (u7_mem_b0_b_106 ), .B (n_3792), .S0 (n_7493), .Y(n_9399));
MX2X1 g34090(.A (u7_mem_b0_b_105 ), .B (n_3645), .S0 (n_7493), .Y(n_8748));
MX2X1 g34097(.A (u7_mem_b0_b_111 ), .B (n_3568), .S0 (n_7493), .Y(n_8740));
MX2X1 g34096(.A (u7_mem_b0_b_110 ), .B (n_3642), .S0 (n_7493), .Y(n_8742));
MX2X1 g34095(.A (u7_mem_b0_b_91 ), .B (n_3566), .S0 (n_7493), .Y(n_8744));
MX2X1 g34094(.A (u7_mem_b0_b_109 ), .B (n_2635), .S0 (n_7493), .Y(n_9398));
MX2X1 g37293(.A (u11_mem_b1_b_145 ), .B (n_5307), .S0 (n_6502), .Y(n_5319));
NAND2X1 g39560(.A (u6_mem_b2_b_35 ), .B (n_2285), .Y (n_1810));
XOR2X1 g40439(.A (n_6316), .B (n_1924), .Y (n_4795));
MX2X1 g40432(.A (crac_din_704), .B (in_slt_843), .S0 (n_1036), .Y(n_1192));
INVX1 g35410(.A (in_valid_s_b0_b ), .Y (n_7389));
INVX1 g35412(.A (n_7356), .Y (n_7357));
INVX1 g35414(.A (in_valid_s_b1_b ), .Y (n_7356));
INVX4 g40455(.A (wb_din_674), .Y (n_2755));
INVX1 g35416(.A (n_7477), .Y (n_7388));
INVX1 g35417(.A (in_valid_s_b2_b ), .Y (n_7477));
AND2X1 g35419(.A (n_5450), .B (u2_sync_resume), .Y (n_6053));
INVX1 g42084(.A (u11_mem_b3_b_72 ), .Y (n_6023));
NAND2X1 g39561(.A (u6_mem_b2_b_51 ), .B (n_3423), .Y (n_3094));
NOR2X1 g39413(.A (n_3453), .B (n_2720), .Y (n_3198));
INVX2 g40476(.A (wb_din_691), .Y (n_2748));
NAND2X1 g39562(.A (u6_mem_b1_b_82 ), .B (n_4253), .Y (n_4167));
INVX2 g32828(.A (n_9737), .Y (n_10303));
INVX4 g32829(.A (n_10073), .Y (n_9737));
MX2X1 g40430(.A (crac_din), .B (in_slt_830), .S0 (n_1036), .Y(n_1074));
INVX4 g32825(.A (n_9737), .Y (n_10267));
NAND2X1 g36949(.A (n_2526), .B (n_1612), .Y (n_4809));
NAND2X1 g39563(.A (u7_mem_b2_b_41 ), .B (n_12641), .Y (n_3093));
INVX1 g42101(.A (oc5_int_set_718), .Y (n_525));
NAND2X1 g52(.A (n_6174), .B (n_12115), .Y (n_12667));
NAND2X1 g51(.A (n_12531), .B (n_6246), .Y (n_11923));
MX2X1 g40431(.A (crac_din_703), .B (in_slt_842), .S0 (n_1036), .Y(n_1193));
NAND2X1 g36948(.A (n_1621), .B (n_1617), .Y (n_4016));
INVX1 g39564(.A (n_4755), .Y (n_3092));
NOR2X1 g40061(.A (n_1147), .B (n_2794), .Y (n_2796));
NOR2X1 g40060(.A (n_2744), .B (n_2182), .Y (n_1805));
NOR2X1 g40063(.A (n_2705), .B (n_2792), .Y (n_2793));
NOR2X1 g40065(.A (n_2729), .B (n_1985), .Y (n_2164));
NOR2X1 g40064(.A (n_1226), .B (n_2790), .Y (n_2791));
NOR2X1 g40066(.A (n_2081), .B (n_2702), .Y (n_2162));
NOR2X1 g40069(.A (n_2788), .B (n_2804), .Y (n_2789));
NOR2X1 g40068(.A (n_2470), .B (n_2818), .Y (n_2161));
AOI21X1 g38399(.A0 (u7_mem_b1_b_64 ), .A1 (n_5069), .B0 (n_2694), .Y(n_4951));
NAND2X1 g39565(.A (in_slt_409), .B (n_2368), .Y (n_4755));
AOI21X1 g38394(.A0 (u8_mem_b2_b_40 ), .A1 (n_4499), .B0 (n_1966), .Y(n_4344));
AOI21X1 g38395(.A0 (u3_mem_b2_b_53 ), .A1 (n_4519), .B0 (n_2084), .Y(n_4343));
AOI21X1 g38396(.A0 (u3_mem_b3_b_152 ), .A1 (n_5133), .B0 (n_3338), .Y(n_4953));
AOI21X1 g38397(.A0 (u7_mem_b3_b_139 ), .A1 (n_4961), .B0 (n_3198), .Y(n_4952));
AOI21X1 g38390(.A0 (u3_mem_b3_b_135 ), .A1 (n_5138), .B0 (n_3478), .Y(n_4955));
AOI21X1 g38391(.A0 (u3_mem_b2_b_51 ), .A1 (n_4519), .B0 (n_2003), .Y(n_4345));
AOI21X1 g38392(.A0 (u8_mem_b3_b_126 ), .A1 (n_3879), .B0 (n_1502), .Y(n_3856));
AOI21X1 g38393(.A0 (u3_mem_b3_b_125 ), .A1 (n_5133), .B0 (n_3391), .Y(n_4954));
XOR2X1 g40437(.A (u11_rp_b1_b ), .B (n_853), .Y (n_1438));
NAND2X1 g39566(.A (u6_mem_b2_b_37 ), .B (n_3474), .Y (n_3091));
NOR2X1 g39567(.A (n_3089), .B (n_2691), .Y (n_3090));
MX2X1 g40435(.A (crac_din_701), .B (in_slt_840), .S0 (n_1036), .Y(n_1031));
NAND2X1 g36672(.A (n_5253), .B (n_2578), .Y (n_5763));
AOI21X1 g37250(.A0 (n_5357), .A1 (n_6594), .B0 (n_3957), .Y (n_5358));
MX2X1 g37251(.A (u10_mem_b1_b_143 ), .B (n_5355), .S0 (n_6475), .Y(n_5356));
AOI21X1 g37253(.A0 (n_5510), .A1 (n_6594), .B0 (n_4658), .Y (n_5511));
AOI21X1 g37254(.A0 (n_5508), .A1 (n_6649), .B0 (n_4643), .Y (n_5509));
AOI21X1 g37256(.A0 (n_5504), .A1 (n_6594), .B0 (n_4655), .Y (n_5505));
AOI21X1 g37257(.A0 (n_5350), .A1 (n_5371), .B0 (n_3953), .Y (n_5351));
AOI21X1 g37258(.A0 (n_5502), .A1 (n_6649), .B0 (n_4640), .Y (n_5503));
AOI21X1 g37259(.A0 (n_5500), .A1 (n_6649), .B0 (n_4652), .Y (n_5501));
AOI21X1 g37704(.A0 (n_256), .A1 (n_2553), .B0 (n_2307), .Y (n_3925));
AOI22X1 g37705(.A0 (n_2558), .A1 (n_337), .B0 (n_5575), .B1 (n_1316),.Y (n_1248));
AOI21X1 g37702(.A0 (n_5577), .A1 (n_1316), .B0 (n_2341), .Y (n_3927));
AOI22X1 g37703(.A0 (n_6548), .A1 (n_1643), .B0 (n_6625), .B1(n_1831), .Y (n_1689));
AOI22X1 g37700(.A0 (n_2558), .A1 (n_314), .B0 (n_1690), .B1 (n_2544),.Y (n_1691));
OAI21X1 g30967(.A0 (n_4788), .A1 (n_10747), .B0 (n_10057), .Y(n_10746));
NAND2X1 g41229(.A (n_601), .B (n_600), .Y (n_602));
NAND2X1 g33018(.A (n_414), .B (n_9882), .Y (n_9884));
OAI21X1 g33019(.A0 (n_753), .A1 (u15_rdd2), .B0 (n_9882), .Y(n_9883));
OAI21X1 g33016(.A0 (n_7260), .A1 (n_7096), .B0 (n_12609), .Y(n_9798));
OAI21X1 g33017(.A0 (n_7258), .A1 (n_7116), .B0 (n_12609), .Y(n_9797));
OAI21X1 g33015(.A0 (n_7262), .A1 (n_7047), .B0 (n_12609), .Y(n_12815));
OAI21X1 g33013(.A0 (n_7126), .A1 (n_7099), .B0 (n_12609), .Y(n_12811));
AOI21X1 g33010(.A0 (crac_wr), .A1 (n_9710), .B0 (u13_ints_r_b1_b ), .Y(n_9803));
OAI21X1 g33011(.A0 (n_7279), .A1 (n_7105), .B0 (n_9885), .Y(n_12008));
NAND2X1 g39431(.A (u10_din_tmp_50), .B (n_2302), .Y (n_2303));
AOI21X1 g35603(.A0 (n_5904), .A1 (n_6117), .B0 (n_12604), .Y(n_7260));
NOR2X1 g39436(.A (n_3486), .B (n_2790), .Y (n_3185));
NAND2X1 g39437(.A (u3_mem_b2_b_56 ), .B (n_3330), .Y (n_3184));
NAND2X1 g31708(.A (n_232), .B (n_10081), .Y (n_9983));
NAND2X1 g31709(.A (n_1684), .B (n_10065), .Y (n_9982));
NAND2X1 g39434(.A (n_12679), .B (u5_mem_b0_b_110 ), .Y (n_3186));
NAND2X1 g40939(.A (n_121), .B (n_4074), .Y (n_1160));
NAND2X1 g40938(.A (n_703), .B (u2_to_cnt_b5_b ), .Y (n_704));
NAND2X1 g31701(.A (n_188), .B (n_10385), .Y (n_10362));
NAND2X1 g31702(.A (n_125), .B (n_10376), .Y (n_10361));
NAND2X1 g31703(.A (n_190), .B (n_10376), .Y (n_10360));
NAND2X1 g31704(.A (n_90), .B (n_10010), .Y (n_9986));
NAND2X1 g31705(.A (n_122), .B (n_10376), .Y (n_10359));
NAND2X1 g31706(.A (n_249), .B (n_10010), .Y (n_9985));
NAND2X1 g31707(.A (n_87), .B (n_10010), .Y (n_9984));
AOI21X1 g38298(.A0 (u5_mem_b1_b_65 ), .A1 (n_5048), .B0 (n_2758), .Y(n_5013));
AOI21X1 g35602(.A0 (n_6140), .A1 (n_5929), .B0 (n_12604), .Y(n_7262));
INVX1 g41089(.A (n_832), .Y (n_1042));
MX2X1 g36143(.A (n_6857), .B (n_6891), .S0 (n_6856), .Y (n_6858));
NAND2X1 g39204(.A (u4_mem_b1_b_64 ), .B (n_12252), .Y (n_11667));
INVX4 g41085(.A (n_1042), .Y (n_6475));
NAND2X1 g34602(.A (u6_mem_b1_b_72 ), .B (n_7758), .Y (n_7827));
INVX1 g42164(.A (u10_mem_b2_b_88 ), .Y (n_6028));
OAI21X1 g33923(.A0 (n_4870), .A1 (n_8911), .B0 (n_7600), .Y (n_8917));
AOI22X1 g37857(.A0 (n_1756), .A1 (n_6347), .B0 (n_6530), .B1(n_1575), .Y (n_1570));
OAI21X1 g33920(.A0 (n_4397), .A1 (n_8933), .B0 (n_7949), .Y (n_8921));
OAI21X1 g33921(.A0 (n_4281), .A1 (n_8891), .B0 (n_7602), .Y (n_8920));
OAI21X1 g33926(.A0 (n_4869), .A1 (n_8911), .B0 (n_7597), .Y (n_8912));
OAI21X1 g33927(.A0 (n_4290), .A1 (n_8930), .B0 (n_7564), .Y (n_8910));
NAND2X1 g36312(.A (n_5893), .B (n_2567), .Y (n_5939));
OAI21X1 g33924(.A0 (n_4280), .A1 (n_8438), .B0 (n_7599), .Y (n_8916));
NAND2X1 g36313(.A (n_5800), .B (n_2567), .Y (n_5938));
OAI21X1 g33925(.A0 (n_4382), .A1 (n_8438), .B0 (n_7598), .Y (n_8914));
INVX1 g42754(.A (u11_mem_b0_b_167 ), .Y (n_334));
INVX1 g42757(.A (u11_mem_b1_b_123 ), .Y (n_6545));
INVX1 g42756(.A (oc0_int_set_707), .Y (n_616));
OAI21X1 g33928(.A0 (n_4868), .A1 (n_8911), .B0 (n_7957), .Y (n_8908));
INVX1 g42753(.A (n_5588), .Y (n_564));
AOI21X1 g35627(.A0 (n_6298), .A1 (n_6122), .B0 (n_12640), .Y(n_7239));
OAI21X1 g33579(.A0 (n_5095), .A1 (n_9346), .B0 (n_7974), .Y (n_9348));
OAI21X1 g33929(.A0 (n_4279), .A1 (n_8930), .B0 (n_7595), .Y (n_8907));
AOI21X1 g35623(.A0 (n_5916), .A1 (n_5759), .B0 (n_7212), .Y (n_7124));
AOI21X1 g35622(.A0 (n_6145), .A1 (n_6283), .B0 (n_7214), .Y (n_7244));
AOI21X1 g35621(.A0 (n_5917), .A1 (n_6104), .B0 (n_7256), .Y (n_7245));
AOI21X1 g35620(.A0 (n_5918), .A1 (n_6105), .B0 (n_7256), .Y (n_7246));
AOI21X1 g35629(.A0 (n_6297), .A1 (n_6119), .B0 (n_12640), .Y(n_7236));
INVX4 g40668(.A (wb_din_676), .Y (n_2786));
NOR2X1 g40232(.A (n_2470), .B (n_2864), .Y (n_2471));
INVX1 g42163(.A (oc2_cfg_986), .Y (n_242));
INVX4 g42287(.A (u6_rp_b0_b ), .Y (n_6821));
MX2X1 g31216(.A (n_6440), .B (n_6439), .S0 (n_10513), .Y (n_10498));
OAI21X1 g33792(.A0 (n_5063), .A1 (n_9080), .B0 (n_7735), .Y (n_9082));
OAI21X1 g33795(.A0 (n_5101), .A1 (n_9077), .B0 (n_7732), .Y (n_9078));
INVX1 g42289(.A (u9_mem_b3_b_57 ), .Y (n_6919));
INVX1 g42579(.A (u11_mem_b0_b_179 ), .Y (n_1585));
NAND2X1 g34251(.A (u8_mem_b3_b_143 ), .B (n_7976), .Y (n_8151));
OAI21X1 g33570(.A0 (n_4407), .A1 (n_8318), .B0 (n_7987), .Y (n_8266));
INVX1 g42571(.A (u11_mem_b3_b_74 ), .Y (n_5580));
INVX1 g42570(.A (u11_mem_b3_b_73 ), .Y (n_6026));
INVX1 g42575(.A (u10_mem_b3_b_58 ), .Y (n_6578));
OAI21X1 g33573(.A0 (n_5105), .A1 (n_8318), .B0 (n_7983), .Y (n_8262));
NAND2X1 g39700(.A (u4_mem_b1_b_69 ), .B (n_12250), .Y (n_11647));
NOR2X1 g39701(.A (n_3117), .B (n_3008), .Y (n_3010));
NOR2X1 g39702(.A (n_2763), .B (n_1488), .Y (n_1476));
NAND2X1 g34252(.A (u8_mem_b3_b_144 ), .B (n_7976), .Y (n_8150));
NAND2X1 g35443(.A (n_5276), .B (n_7113), .Y (n_7338));
INVX1 g39705(.A (n_4761), .Y (n_2886));
NAND2X1 g39706(.A (n_2302), .B (in_slt_432), .Y (n_4761));
NAND2X1 g39708(.A (in_slt_401), .B (n_2368), .Y (n_2259));
OAI21X1 g33575(.A0 (n_5103), .A1 (n_9349), .B0 (n_7980), .Y (n_8260));
OAI21X1 g33574(.A0 (n_5104), .A1 (n_8318), .B0 (n_7981), .Y (n_8261));
MX2X1 g31332(.A (n_6348), .B (n_6347), .S0 (n_10537), .Y (n_10417));
NOR2X1 g36828(.A (n_5736), .B (n_5371), .Y (n_5570));
NAND2X1 g34257(.A (u7_mem_b2_b_57 ), .B (n_7651), .Y (n_8145));
AOI21X1 g40234(.A0 (ic0_cfg_1024), .A1 (n_221), .B0(u14_u6_full_empty_r), .Y (n_843));
NAND4X1 g36824(.A (n_12799), .B (n_3192), .C (n_12800), .D (n_1338),.Y (n_5859));
NAND2X1 g36825(.A (n_1657), .B (n_2554), .Y (n_4822));
INVX1 g36826(.A (n_6266), .Y (n_5727));
OAI21X1 g33576(.A0 (n_5099), .A1 (n_9349), .B0 (n_7979), .Y (n_8259));
NAND2X1 g36820(.A (n_1840), .B (n_2555), .Y (n_4823));
NAND4X1 g36822(.A (n_11662), .B (n_11663), .C (n_2644), .D (n_3533),.Y (n_6246));
INVX1 g36823(.A (n_5859), .Y (n_5571));
NOR2X1 g35442(.A (n_7022), .B (n_3431), .Y (n_7023));
NOR2X1 g40830(.A (n_4734), .B (n_936), .Y (n_8843));
NAND2X1 g40831(.A (n_4734), .B (n_936), .Y (n_7524));
NOR2X1 g35441(.A (n_7025), .B (n_1216), .Y (n_7024));
NAND2X1 g39403(.A (u5_mem_b2_b_59 ), .B (n_12823), .Y (n_1624));
NAND2X1 g36429(.A (n_6794), .B (n_12531), .Y (n_6809));
NAND2X1 g37951(.A (n_2379), .B (n_3184), .Y (n_5188));
NAND2X1 g37953(.A (n_1811), .B (n_3495), .Y (n_5187));
NAND2X1 g37957(.A (n_2888), .B (n_3840), .Y (n_5183));
NAND2X1 g35447(.A (n_7300), .B (n_6694), .Y (n_7454));
NAND2X1 g37956(.A (n_2871), .B (n_2984), .Y (n_5184));
NAND2X1 g37955(.A (n_2464), .B (n_3122), .Y (n_5185));
NAND2X1 g37954(.A (n_3045), .B (n_3004), .Y (n_5186));
OAI21X1 g33830(.A0 (n_4893), .A1 (n_8981), .B0 (n_7692), .Y (n_9033));
OAI21X1 g33831(.A0 (n_5009), .A1 (n_9055), .B0 (n_7906), .Y (n_9031));
OAI21X1 g33832(.A0 (n_4892), .A1 (n_8948), .B0 (n_7691), .Y (n_9030));
OAI21X1 g33833(.A0 (n_5117), .A1 (n_9034), .B0 (n_7690), .Y (n_9029));
OAI21X1 g33834(.A0 (n_4951), .A1 (n_9034), .B0 (n_7689), .Y (n_9028));
OAI21X1 g33835(.A0 (n_5070), .A1 (n_9043), .B0 (n_7688), .Y (n_9026));
NAND2X1 g34288(.A (u3_mem_b2_b_32 ), .B (n_8141), .Y (n_8112));
NAND2X1 g34289(.A (u3_mem_b2_b_33 ), .B (n_8141), .Y (n_8110));
NAND2X1 g34286(.A (u3_mem_b2_b_59 ), .B (n_8101), .Y (n_8114));
NAND2X1 g34287(.A (u3_mem_b2_b_31 ), .B (n_8101), .Y (n_8113));
NAND2X1 g34284(.A (u3_mem_b2_b_30 ), .B (n_8101), .Y (n_8116));
NAND2X1 g34285(.A (u3_mem_b2_b_58 ), .B (n_8141), .Y (n_8115));
NAND2X1 g34282(.A (u8_mem_b3_b ), .B (n_7976), .Y (n_8118));
NAND2X1 g34283(.A (u3_mem_b2_b_57 ), .B (n_8141), .Y (n_8117));
NAND2X1 g34280(.A (u3_mem_b2_b_55 ), .B (n_8141), .Y (n_8120));
NAND2X1 g34281(.A (u3_mem_b2_b_56 ), .B (n_8141), .Y (n_8119));
NAND2X1 g36423(.A (n_5805), .B (n_6152), .Y (n_5897));
AOI21X1 g38086(.A0 (u8_mem_b2_b_32 ), .A1 (n_4499), .B0 (n_2165), .Y(n_4487));
NAND2X1 g36424(.A (n_5895), .B (n_6259), .Y (n_5896));
AOI21X1 g38087(.A0 (u3_mem_b2_b_46 ), .A1 (n_4533), .B0 (n_1983), .Y(n_4486));
NOR2X1 g39653(.A (n_3453), .B (n_2744), .Y (n_3032));
NAND2X1 g36425(.A (n_5893), .B (n_6259), .Y (n_5894));
AOI21X1 g38088(.A0 (u8_mem_b3_b_130 ), .A1 (n_3879), .B0 (n_1470), .Y(n_3877));
NOR2X1 g36426(.A (n_838), .B (n_6057), .Y (n_5892));
AOI21X1 g38089(.A0 (u8_mem_b2_b_31 ), .A1 (n_4491), .B0 (n_2149), .Y(n_4485));
NAND2X1 g35445(.A (n_7386), .B (n_7012), .Y (n_7456));
MX2X1 g36135(.A (n_6402), .B (n_6618), .S0 (n_6856), .Y (n_6403));
NOR2X1 g37506(.A (n_4759), .B (n_6594), .Y (n_3957));
NAND2X1 g37507(.A (n_5480), .B (n_3092), .Y (n_4659));
MX2X1 g38732(.A (u6_mem_b0_b_110 ), .B (wb_din_680), .S0 (n_3632), .Y(n_3609));
NAND2X1 g39406(.A (n_3259), .B (u5_mem_b0_b_109 ), .Y (n_3205));
NOR2X1 g37503(.A (n_5287), .B (n_6594), .Y (n_4661));
NOR2X1 g40006(.A (n_2216), .B (n_2794), .Y (n_2204));
NOR2X1 g40003(.A (n_2169), .B (n_2804), .Y (n_2206));
INVX4 g41129(.A (n_1045), .Y (n_4783));
AND2X1 g37056(.A (n_1553), .B (n_1281), .Y (n_1282));
INVX4 g45590_dup(.A (n_12244), .Y (n_12840));
AND2X1 g40978(.A (n_689), .B (u9_wp_b2_b ), .Y (n_930));
NAND2X1 g32619(.A (n_853), .B (n_9631), .Y (n_9835));
NOR2X1 g32618(.A (n_8476), .B (n_5825), .Y (n_9464));
NOR2X1 g32617(.A (n_8477), .B (n_11086), .Y (n_9465));
NOR2X1 g32616(.A (n_8480), .B (n_5839), .Y (n_9466));
NOR2X1 g32615(.A (n_8478), .B (n_10994), .Y (n_9467));
NOR2X1 g32613(.A (n_8481), .B (n_11030), .Y (n_9469));
NAND2X1 g32612(.A (n_9448), .B (oc5_int_set_718), .Y (n_9573));
NAND2X1 g32611(.A (n_9449), .B (oc4_int_set_716), .Y (n_9574));
NAND2X1 g32610(.A (n_9450), .B (oc3_int_set_714), .Y (n_9575));
NAND4X1 g37067(.A (n_11721), .B (n_11722), .C (n_3341), .D (n_2397),.Y (n_6194));
INVX1 g37066(.A (n_6194), .Y (n_5683));
NAND4X1 g37065(.A (n_3278), .B (n_3000), .C (n_3289), .D (n_1323), .Y(n_6163));
INVX1 g37064(.A (n_6163), .Y (n_5684));
OAI21X1 g33612(.A0 (n_5038), .A1 (n_9307), .B0 (n_7933), .Y (n_9306));
MX2X1 g38701(.A (u6_mem_b0_b_94 ), .B (wb_din_664), .S0 (n_3632), .Y(n_3648));
MX2X1 g38700(.A (u8_mem_b0_b_98 ), .B (wb_din_668), .S0 (n_3826), .Y(n_3649));
NAND4X1 g37069(.A (n_11461), .B (n_11462), .C (n_2237), .D (n_2387),.Y (n_5809));
INVX1 g37068(.A (n_5809), .Y (n_5537));
OAI21X1 g36622(.A0 (n_4568), .A1 (n_5463), .B0 (n_6134), .Y (n_6135));
OAI21X1 g36623(.A0 (n_4611), .A1 (n_5163), .B0 (n_6152), .Y (n_5794));
OAI21X1 g36620(.A0 (n_4569), .A1 (n_5196), .B0 (n_6131), .Y (n_6137));
OAI21X1 g36621(.A0 (n_4632), .A1 (n_5454), .B0 (n_6134), .Y (n_6136));
OAI21X1 g36626(.A0 (n_5165), .A1 (n_5164), .B0 (n_6152), .Y (n_5793));
NAND2X1 g36627(.A (n_5278), .B (n_3982), .Y (n_5791));
OAI21X1 g36624(.A0 (n_4586), .A1 (n_5212), .B0 (n_6134), .Y (n_6133));
OAI21X1 g36625(.A0 (n_4603), .A1 (n_5224), .B0 (n_6131), .Y (n_6132));
AOI21X1 g36628(.A0 (n_5591), .A1 (ic2_cfg_1044), .B0 (n_4681), .Y(n_5592));
INVX1 g43047(.A (n_8199), .Y (n_804));
OAI22X1 g30750(.A0 (n_11097), .A1 (n_5536), .B0 (out_slt9), .B1(n_11096), .Y (n_11102));
OAI22X1 g30751(.A0 (n_11100), .A1 (n_5676), .B0 (n_11099), .B1(out_slt_65), .Y (n_11101));
OAI22X1 g30752(.A0 (n_11097), .A1 (n_5670), .B0 (n_11096), .B1(out_slt_160), .Y (n_11098));
OAI21X1 g37391(.A0 (u10_mem_b0_b_171 ), .A1 (n_6341), .B0 (n_5235), .Y(n_5662));
OAI21X1 g37390(.A0 (u11_mem_b0_b_170 ), .A1 (n_6359), .B0 (n_5242), .Y(n_5664));
OAI21X1 g37393(.A0 (u11_mem_b0_b_180 ), .A1 (n_6359), .B0 (n_5244), .Y(n_5659));
OAI21X1 g37392(.A0 (u11_mem_b0_b_176 ), .A1 (n_6359), .B0 (n_5236), .Y(n_5660));
OAI21X1 g37395(.A0 (u11_mem_b0_b_169 ), .A1 (n_5656), .B0 (n_5245), .Y(n_5657));
OAI21X1 g37394(.A0 (u11_mem_b0_b_178 ), .A1 (n_5656), .B0 (n_5233), .Y(n_5658));
OAI21X1 g37397(.A0 (u11_mem_b0_b_172 ), .A1 (n_6359), .B0 (n_5241), .Y(n_5653));
OAI21X1 g37396(.A0 (u11_mem_b0_b_171 ), .A1 (n_6359), .B0 (n_5246), .Y(n_5655));
OAI21X1 g37399(.A0 (u10_mem_b0_b_170 ), .A1 (n_6341), .B0 (n_4642), .Y(n_5472));
OAI21X1 g37398(.A0 (u11_mem_b0_b_174 ), .A1 (n_6359), .B0 (n_5238), .Y(n_5651));
AOI21X1 g38569(.A0 (u8_mem_b2_b_46 ), .A1 (n_4491), .B0 (n_2056), .Y(n_4272));
AOI21X1 g38568(.A0 (u3_mem_b1_b_60 ), .A1 (n_5148), .B0 (n_2814), .Y(n_4863));
AOI21X1 g35567(.A0 (n_6309), .A1 (n_6136), .B0 (n_12145), .Y(n_7277));
NOR2X1 g39525(.A (n_3117), .B (n_2748), .Y (n_3118));
NOR2X1 g39526(.A (n_4996), .B (n_2804), .Y (n_3116));
NOR2X1 g39241(.A (n_2707), .B (n_1488), .Y (n_1490));
NAND2X1 g41655(.A (u10_rp_b1_b ), .B (u10_wp_b2_b ), .Y (n_480));
AND2X1 g41654(.A (n_693), .B (n_942), .Y (n_9659));
MX2X1 g31393(.A (u10_din_tmp_56), .B (in_slt_437), .S0 (n_9860), .Y(n_9854));
MX2X1 g31392(.A (u10_din_tmp_55), .B (in_slt_436), .S0 (n_9860), .Y(n_9855));
MX2X1 g31391(.A (u10_din_tmp_54), .B (in_slt_435), .S0 (n_9860), .Y(n_9856));
MX2X1 g31390(.A (u10_din_tmp_53), .B (in_slt_434), .S0 (n_9860), .Y(n_9857));
XOR2X1 g31397(.A (n_1012), .B (n_10329), .Y (n_10095));
AOI21X1 g31396(.A0 (n_12339), .A1 (n_1096), .B0 (n_10068), .Y(n_10404));
AOI21X1 g31395(.A0 (n_11893), .A1 (n_757), .B0 (n_10085), .Y(n_10405));
MX2X1 g31394(.A (u10_din_tmp_42), .B (in_slt_423), .S0 (n_9860), .Y(n_9853));
AOI21X1 g31399(.A0 (n_11891), .A1 (n_11586), .B0 (n_9990), .Y(n_10403));
XOR2X1 g31398(.A (n_641), .B (n_10327), .Y (n_10094));
NAND2X1 g37935(.A (n_2911), .B (n_2856), .Y (n_5195));
NAND2X1 g39240(.A (u7_mem_b1_b_61 ), .B (n_4225), .Y (n_4210));
NAND2X1 g37936(.A (n_4222), .B (n_3044), .Y (n_5453));
NAND2X1 g37931(.A (n_4177), .B (n_3516), .Y (n_5454));
NAND2X1 g37930(.A (n_1522), .B (n_4116), .Y (n_5455));
AOI22X1 g37933(.A0 (u10_din_tmp_45), .A1 (n_3339), .B0 (n_3911), .B1(in_slt_424), .Y (n_4557));
AOI22X1 g37932(.A0 (n_385), .A1 (n_1835), .B0 (n_5365), .B1 (n_1760),.Y (n_1858));
NOR2X1 g39023(.A (n_3486), .B (n_3008), .Y (n_3506));
AOI22X1 g37939(.A0 (n_343), .A1 (n_1835), .B0 (n_5350), .B1 (n_1760),.Y (n_2505));
AOI22X1 g37938(.A0 (u10_din_tmp_48), .A1 (n_3339), .B0 (n_3911), .B1(in_slt_427), .Y (n_4555));
INVX1 g33225(.A (o6_empty), .Y (n_9538));
NOR2X1 g41144(.A (n_8188), .B (n_921), .Y (n_9697));
INVX1 g33227(.A (o7_empty), .Y (n_9536));
INVX1 g41410(.A (n_847), .Y (n_1130));
INVX1 g33221(.A (o3_empty), .Y (n_9543));
NAND2X1 g41416(.A (u11_rp_b1_b ), .B (u11_rp_b0_b ), .Y (n_736));
INVX1 g33223(.A (o4_empty), .Y (n_9541));
INVX1 g41142(.A (n_781), .Y (n_1149));
NAND2X1 g41419(.A (u9_rp_b1_b ), .B (u9_rp_b0_b ), .Y (n_737));
INVX1 g33229(.A (o8_empty), .Y (n_9534));
INVX4 g41148(.A (n_1148), .Y (n_2325));
INVX1 g42140(.A (u11_mem_b3_b_66 ), .Y (n_6428));
NAND3X1 g34709(.A (n_4734), .B (n_4736), .C (n_864), .Y (n_1886));
OR2X1 g34708(.A (i4_status), .B (n_7380), .Y (n_7381));
NAND3X1 g34879(.A (n_7499), .B (n_1450), .C (n_991), .Y (n_8677));
NOR2X1 g34878(.A (n_7367), .B (n_4802), .Y (n_7513));
NAND2X1 g34875(.A (u3_mem_b1_b_86 ), .B (n_8141), .Y (n_7559));
NAND2X1 g34874(.A (u8_mem_b2_b_58 ), .B (n_7976), .Y (n_7560));
NAND3X1 g34877(.A (n_7490), .B (n_1454), .C (n_8182), .Y (n_8678));
NAND2X1 g34876(.A (u8_mem_b2_b_31 ), .B (n_7976), .Y (n_7558));
NAND2X1 g34707(.A (n_7382), .B (n_7380), .Y (n_7529));
NAND2X1 g34870(.A (u8_mem_b1_b_88 ), .B (n_7976), .Y (n_7564));
NAND2X1 g34873(.A (u8_mem_b2_b_30 ), .B (n_7976), .Y (n_7561));
NAND2X1 g34872(.A (u3_mem_b1_b_85 ), .B (n_8101), .Y (n_7562));
NAND2X1 g31579(.A (n_2556), .B (n_10010), .Y (n_10078));
NAND2X1 g31578(.A (n_39), .B (n_10010), .Y (n_10079));
NAND2X1 g31577(.A (n_98), .B (n_10081), .Y (n_10080));
NAND2X1 g31576(.A (n_256), .B (n_10081), .Y (n_10082));
NAND2X1 g31575(.A (n_1690), .B (n_10081), .Y (n_10084));
NOR2X1 g31574(.A (n_11894), .B (n_757), .Y (n_10085));
NAND3X1 g31573(.A (u11_wp_b0_b ), .B (n_11772), .C (n_9631), .Y(n_10086));
NAND2X1 g31572(.A (n_4797), .B (n_11126), .Y (n_11509));
NAND2X1 g31571(.A (n_4799), .B (n_11131), .Y (n_11511));
NAND2X1 g31570(.A (n_4795), .B (n_11136), .Y (n_10397));
NOR2X1 g39937(.A (n_3486), .B (n_2864), .Y (n_2865));
NAND2X1 g39936(.A (n_11789), .B (u8_mem_b0_b_93 ), .Y (n_12039));
NAND2X1 g39935(.A (n_3339), .B (in_slt_436), .Y (n_5330));
INVX1 g39934(.A (n_5330), .Y (n_4108));
NAND2X1 g39933(.A (u4_mem_b2_b_35 ), .B (n_12087), .Y (n_2233));
NAND2X1 g39932(.A (u4_mem_b1_b_84 ), .B (n_12250), .Y (n_4109));
NAND2X1 g39931(.A (u8_mem_b1_b_84 ), .B (n_12291), .Y (n_2867));
NAND2X1 g39930(.A (n_11798), .B (u8_mem_b0_b_109 ), .Y (n_2868));
OR2X1 g39939(.A (n_7214), .B (n_6316), .Y (n_2232));
NAND2X1 g39938(.A (u8_mem_b2_b_49 ), .B (n_3441), .Y (n_2863));
MX2X1 g37219(.A (u9_mem_b1_b_139 ), .B (n_4747), .S0 (n_5730), .Y(n_4790));
NAND2X1 g38881(.A (u7_mem_b3_b_136 ), .B (n_1538), .Y (n_1533));
NAND2X1 g38882(.A (u6_mem_b3_b ), .B (n_2419), .Y (n_2431));
AOI21X1 g38244(.A0 (u6_mem_b3_b_150 ), .A1 (n_5100), .B0 (n_3235), .Y(n_5061));
NAND2X1 g38883(.A (u5_mem_b3_b_150 ), .B (n_3543), .Y (n_3536));
NAND2X1 g38884(.A (u6_mem_b3_b_127 ), .B (n_2419), .Y (n_1869));
NAND2X1 g38885(.A (u6_mem_b3_b_143 ), .B (n_2465), .Y (n_2429));
NAND2X1 g38834(.A (u3_mem_b3_b_128 ), .B (n_1517), .Y (n_1323));
NAND2X1 g38886(.A (u6_mem_b3_b_129 ), .B (n_2419), .Y (n_2428));
NAND2X1 g38887(.A (u5_mem_b3_b_131 ), .B (n_1543), .Y (n_1340));
NOR2X1 g39247(.A (n_2765), .B (n_1488), .Y (n_1489));
AOI22X1 g30118(.A0 (n_9583), .A1 (n_9611), .B0 (n_752), .B1 (n_9503),.Y (n_9755));
AOI22X1 g30119(.A0 (n_9643), .A1 (n_9656), .B0 (n_683), .B1 (n_9560),.Y (n_9837));
AOI21X1 g35568(.A0 (n_5897), .A1 (n_6324), .B0 (n_7120), .Y (n_7276));
AOI21X1 g35472(.A0 (i4_dout_616), .A1 (n_7468), .B0 (n_7135), .Y(n_7332));
AOI21X1 g35473(.A0 (i3_dout_579), .A1 (n_6700), .B0 (n_7134), .Y(n_7331));
AOI21X1 g35470(.A0 (i3_dout_583), .A1 (n_6700), .B0 (n_7137), .Y(n_7335));
OR2X1 g30111(.A (u13_ints_r_b26_b ), .B (ic2_int_set), .Y (n_9757));
AOI22X1 g30116(.A0 (n_9584), .A1 (n_9614), .B0 (n_672), .B1(n_12847), .Y (n_9756));
AOI22X1 g30117(.A0 (n_9644), .A1 (n_9659), .B0 (n_741), .B1(n_12845), .Y (n_9838));
AOI21X1 g35474(.A0 (u10_rp_b1_b ), .A1 (i4_re), .B0 (n_6707), .Y(n_7150));
NOR2X1 g35475(.A (i3_empty), .B (i3_re), .Y (n_7149));
NAND2X1 g39548(.A (u7_mem_b1_b_72 ), .B (n_11856), .Y (n_4173));
MX2X1 g31290(.A (n_6369), .B (n_6368), .S0 (n_9818), .Y (n_10815));
INVX1 g42691(.A (u10_mem_b3_b_65 ), .Y (n_6000));
NAND2X1 g32842(.A (n_12148), .B (n_12144), .Y (n_10992));
NOR2X1 g32843(.A (n_9626), .B (n_12144), .Y (n_10329));
NAND3X1 g32840(.A (n_9690), .B (n_4680), .C (n_11564), .Y (n_9734));
NAND3X1 g32841(.A (n_9620), .B (n_5250), .C (n_11600), .Y (n_9831));
NOR2X1 g32846(.A (n_12603), .B (n_11491), .Y (n_10327));
NOR2X1 g32844(.A (n_9364), .B (n_10940), .Y (n_9518));
NAND2X1 g32845(.A (n_12607), .B (n_12603), .Y (n_10985));
NAND2X1 g34343(.A (u3_mem_b2_b_50 ), .B (n_8101), .Y (n_8060));
AOI22X1 g45892(.A0 (u6_mem_b2_b_42 ), .A1 (n_2285), .B0 (n_12622), .B1(u6_mem_b3_b_135 ), .Y (n_12623));
INVX1 g42698(.A (u4_wp_b1_b ), .Y (n_444));
NAND2X1 g39546(.A (u4_mem_b2_b_39 ), .B (n_12079), .Y (n_1808));
NAND3X1 g45891(.A (n_12623), .B (n_12624), .C (n_12625), .Y(n_12626));
INVX1 g45362(.A (n_11586), .Y (n_11585));
NAND2X1 g34342(.A (u3_mem_b3_b_144 ), .B (n_8097), .Y (n_8061));
NAND2X1 g40049(.A (n_5048), .B (n_4378), .Y (n_2175));
NOR2X1 g40043(.A (n_1226), .B (n_2772), .Y (n_2807));
NOR2X1 g40042(.A (n_2093), .B (n_2686), .Y (n_2178));
NOR2X1 g40041(.A (n_2470), .B (n_2681), .Y (n_2180));
NOR2X1 g40040(.A (n_2827), .B (n_2767), .Y (n_2808));
NOR2X1 g40047(.A (n_2054), .B (n_2782), .Y (n_2177));
NOR2X1 g40046(.A (n_969), .B (n_930), .Y (n_1209));
NAND2X1 g34341(.A (u8_mem_b2_b_59 ), .B (n_7976), .Y (n_8062));
NOR2X1 g40044(.A (n_941), .B (n_2729), .Y (n_1800));
NAND2X1 g34340(.A (u3_mem_b3_b_145 ), .B (n_8097), .Y (n_8063));
NAND2X1 g39313(.A (u6_mem_b2_b_48 ), .B (n_3423), .Y (n_3283));
INVX2 g40554(.A (wb_din_669), .Y (n_2686));
NAND2X1 g34347(.A (n_6691), .B (n_7469), .Y (n_8234));
MX2X1 g40436(.A (crac_din_692), .B (in_slt_831), .S0 (n_1036), .Y(n_1202));
NAND2X1 g34346(.A (u3_mem_b3_b_125 ), .B (n_8101), .Y (n_8057));
AOI22X1 g37728(.A0 (n_9), .A1 (n_2544), .B0 (n_5514), .B1 (n_1316),.Y (n_1683));
AOI22X1 g37729(.A0 (n_3911), .A1 (in_slt_429), .B0 (n_2344), .B1(in_slt_427), .Y (n_2552));
AOI21X1 g37238(.A0 (n_5369), .A1 (n_5371), .B0 (n_3963), .Y (n_5370));
AOI21X1 g37239(.A0 (n_5367), .A1 (n_5371), .B0 (n_3952), .Y (n_5368));
NAND2X1 g34345(.A (u3_mem_b1_b_66 ), .B (n_8141), .Y (n_8058));
INVX1 g35147(.A (n_7402), .Y (n_9043));
MX2X1 g37232(.A (u9_mem_b2_b_115 ), .B (n_4772), .S0 (n_6898), .Y(n_4773));
MX2X1 g37233(.A (u9_mem_b2_b_116 ), .B (n_4769), .S0 (n_6898), .Y(n_4770));
MX2X1 g37230(.A (u9_mem_b2_b_111 ), .B (n_4753), .S0 (n_5732), .Y(n_4775));
MX2X1 g37231(.A (u9_mem_b2_b_113 ), .B (n_4749), .S0 (n_6898), .Y(n_4774));
AOI21X1 g37236(.A0 (n_5374), .A1 (n_5371), .B0 (n_4085), .Y (n_5375));
AOI21X1 g37237(.A0 (n_5372), .A1 (n_5371), .B0 (n_3949), .Y (n_5373));
MX2X1 g37234(.A (u9_mem_b2_b_118 ), .B (n_4767), .S0 (n_6898), .Y(n_4768));
MX2X1 g37235(.A (u10_mem_b1_b_144 ), .B (n_4761), .S0 (n_5407), .Y(n_4766));
OAI21X1 g33038(.A0 (n_12632), .A1 (n_7091), .B0 (n_12161), .Y(n_10209));
OAI21X1 g33039(.A0 (n_12639), .A1 (n_7090), .B0 (n_12161), .Y(n_10207));
OAI21X1 g33030(.A0 (n_7248), .A1 (n_7184), .B0 (n_10518), .Y(n_11956));
OAI21X1 g33031(.A0 (n_7312), .A1 (n_7092), .B0 (n_10518), .Y(n_11958));
OAI21X1 g33032(.A0 (n_7311), .A1 (n_6991), .B0 (n_10518), .Y(n_11996));
OAI21X1 g33033(.A0 (n_7309), .A1 (n_6990), .B0 (n_10518), .Y(n_11960));
OAI21X1 g33034(.A0 (n_7246), .A1 (n_6989), .B0 (n_10518), .Y(n_11962));
OAI21X1 g33035(.A0 (n_7245), .A1 (n_7183), .B0 (n_10518), .Y(n_11976));
OAI21X1 g33036(.A0 (n_7318), .A1 (n_12359), .B0 (n_12149), .Y(n_12000));
OAI21X1 g33037(.A0 (n_7278), .A1 (n_7046), .B0 (n_12149), .Y(n_12010));
NAND2X1 g34344(.A (n_6738), .B (n_7470), .Y (n_8235));
INVX1 g40959(.A (n_1427), .Y (n_2759));
INVX1 g40958(.A (n_1427), .Y (n_2770));
BUFX3 g40951(.A (n_1082), .Y (n_5048));
NOR2X1 g40950(.A (n_8526), .B (n_924), .Y (n_9701));
BUFX3 g40952(.A (n_1082), .Y (n_5037));
INVX1 g40955(.A (n_1427), .Y (n_2773));
INVX2 g40954(.A (n_1427), .Y (n_2784));
INVX2 g40957(.A (n_1082), .Y (n_1427));
INVX1 g40956(.A (n_1427), .Y (n_2827));
NAND2X1 g38956(.A (u3_mem_b3_b_131 ), .B (n_1517), .Y (n_1513));
NAND2X1 g38957(.A (u4_mem_b3_b_128 ), .B (n_12744), .Y (n_4251));
NAND2X1 g38954(.A (u3_mem_b3_b ), .B (n_1517), .Y (n_1514));
NAND2X1 g38952(.A (u3_mem_b3_b_136 ), .B (n_1517), .Y (n_1515));
NAND2X1 g39278(.A (n_12721), .B (u3_mem_b0_b_99 ), .Y (n_12005));
NAND2X1 g34264(.A (u8_mem_b3_b_124 ), .B (n_7976), .Y (n_8137));
NOR2X1 g35814(.A (n_696), .B (n_6752), .Y (n_6746));
INVX1 g42772(.A (u11_rp_b1_b ), .Y (n_5));
NOR2X1 g35815(.A (n_612), .B (n_6752), .Y (n_6672));
NOR2X1 g35816(.A (n_580), .B (n_5440), .Y (n_6747));
INVX1 g42779(.A (u10_mem_b0_b_156 ), .Y (n_6333));
OAI21X1 g36670(.A0 (n_12054), .A1 (n_12055), .B0 (n_784), .Y(n_6116));
NAND3X1 g31762(.A (n_12115), .B (n_12689), .C (n_862), .Y (n_11100));
AOI21X1 g31763(.A0 (n_1500), .A1 (n_4080), .B0 (n_11890), .Y(n_9967));
AOI21X1 g31760(.A0 (n_9672), .A1 (i6_full), .B0 (n_749), .Y(n_10341));
AND2X1 g31761(.A (n_1778), .B (ac97_rst_force), .Y (n_9491));
AOI21X1 g31766(.A0 (n_1122), .A1 (n_7037), .B0 (n_12848), .Y(n_9556));
NAND3X1 g31764(.A (n_6259), .B (n_10483), .C (n_8182), .Y (n_11097));
INVX1 g31765(.A (n_9556), .Y (n_9557));
AOI21X1 g31768(.A0 (n_1127), .A1 (n_7161), .B0 (n_12846), .Y(n_9606));
INVX1 g31769(.A (n_9554), .Y (n_9555));
NOR2X1 g35811(.A (n_677), .B (n_5440), .Y (n_6742));
AOI21X1 g35641(.A0 (n_6290), .A1 (n_5753), .B0 (n_7214), .Y (n_7225));
OAI21X1 g35864(.A0 (n_6081), .A1 (n_11934), .B0 (n_6809), .Y(n_7196));
OAI21X1 g35867(.A0 (n_5725), .A1 (n_11934), .B0 (n_6253), .Y(n_7104));
NAND2X1 g39893(.A (u4_mem_b2_b_52 ), .B (n_12091), .Y (n_2897));
AOI21X1 g35645(.A0 (n_6288), .A1 (n_5796), .B0 (n_7214), .Y (n_7219));
OAI21X1 g35860(.A0 (n_6073), .A1 (n_11934), .B0 (n_6812), .Y(n_7201));
OAI21X1 g35863(.A0 (n_5678), .A1 (n_11934), .B0 (n_6810), .Y(n_7292));
AOI21X1 g35646(.A0 (n_5913), .A1 (n_6093), .B0 (n_7212), .Y (n_7218));
AOI21X1 g35649(.A0 (n_5911), .A1 (n_5748), .B0 (n_7212), .Y (n_7122));
AOI21X1 g35648(.A0 (n_6287), .A1 (n_5749), .B0 (n_7214), .Y (n_7217));
NOR2X1 g35813(.A (n_669), .B (n_6752), .Y (n_6744));
OAI21X1 g35869(.A0 (n_5729), .A1 (n_11934), .B0 (n_6249), .Y(n_7103));
OAI21X1 g35868(.A0 (n_5724), .A1 (n_11934), .B0 (n_6793), .Y(n_7194));
NAND2X1 g39540(.A (n_12839), .B (u4_mem_b0_b_112 ), .Y (n_3104));
NAND2X1 g39541(.A (n_2491), .B (u7_mem_b0_b_93 ), .Y (n_2289));
NAND2X1 g36355(.A (n_5847), .B (n_6821), .Y (n_5921));
NAND2X1 g34266(.A (u8_mem_b3_b_125 ), .B (n_7976), .Y (n_8134));
INVX1 g42479(.A (u10_mem_b3_b_66 ), .Y (n_6601));
INVX1 g42553(.A (u10_mem_b1_b_146 ), .Y (n_215));
INVX1 g42552(.A (u11_mem_b0_b_150 ), .Y (n_6388));
INVX1 g42551(.A (u10_mem_b2_b_100 ), .Y (n_6664));
INVX1 g42550(.A (oc4_cfg_1006), .Y (n_528));
INVX1 g42557(.A (u10_mem_b1_b_133 ), .Y (n_502));
INVX1 g42558(.A (u11_mem_b2_b_112 ), .Y (n_270));
NAND2X1 g9(.A (n_12331), .B (n_12332), .Y (n_12333));
MX2X1 g38757(.A (u3_mem_b0_b_120 ), .B (wb_din_690), .S0 (n_3807), .Y(n_3579));
NAND2X1 g39768(.A (u7_mem_b1_b_69 ), .B (n_4130), .Y (n_4131));
NAND2X1 g39769(.A (u5_mem_b1_b_68 ), .B (n_1035), .Y (n_3194));
INVX1 g39762(.A (n_5304), .Y (n_4133));
INVX1 g39422(.A (n_5296), .Y (n_4193));
NOR2X1 g39092(.A (n_3453), .B (n_2786), .Y (n_3455));
NAND2X1 g39761(.A (u4_mem_b1_b_88 ), .B (n_12267), .Y (n_4134));
NOR2X1 g39094(.A (n_3453), .B (n_2712), .Y (n_3454));
NAND2X1 g39095(.A (u7_mem_b2_b_49 ), .B (n_12654), .Y (n_3452));
NAND2X1 g36353(.A (n_6207), .B (n_12634), .Y (n_6308));
NOR2X1 g39097(.A (n_3117), .B (n_2732), .Y (n_3449));
INVX1 g41902(.A (u11_wp_b0_b ), .Y (n_393));
XOR2X1 g38240(.A (n_95), .B (n_5102), .Y (n_4395));
INVX1 g42302(.A (n_705), .Y (n_6841));
MX2X1 g31186(.A (n_6499), .B (n_6498), .S0 (n_9721), .Y (n_10554));
MX2X1 g31187(.A (n_6493), .B (n_6492), .S0 (n_10513), .Y (n_10552));
MX2X1 g31184(.A (n_5989), .B (n_5988), .S0 (n_10513), .Y (n_10556));
MX2X1 g31185(.A (n_6501), .B (n_6500), .S0 (n_9721), .Y (n_10555));
MX2X1 g31182(.A (n_6504), .B (n_6503), .S0 (n_10513), .Y (n_10558));
MX2X1 g31183(.A (n_5991), .B (n_5990), .S0 (n_9818), .Y (n_10842));
MX2X1 g31180(.A (n_6512), .B (n_6511), .S0 (n_10820), .Y (n_10843));
MX2X1 g31181(.A (n_6508), .B (n_6507), .S0 (n_10513), .Y (n_10559));
NAND2X1 g39306(.A (in_slt_398), .B (n_3415), .Y (n_3291));
NAND2X1 g38830(.A (u5_mem_b3_b_128 ), .B (n_1543), .Y (n_1548));
MX2X1 g31188(.A (n_6491), .B (n_6490), .S0 (n_10513), .Y (n_10551));
MX2X1 g31189(.A (n_6546), .B (n_6545), .S0 (n_10513), .Y (n_10549));
NAND2X1 g34261(.A (u8_mem_b3_b_123 ), .B (n_7976), .Y (n_8140));
MX2X1 g34149(.A (u8_mem_b0_b_117 ), .B (n_3651), .S0 (n_7490), .Y(n_8695));
INVX1 g41908(.A (u7_wp_b0_b ), .Y (n_746));
NAND2X1 g34262(.A (u8_mem_b3_b_151 ), .B (n_7976), .Y (n_8139));
MX2X1 g34118(.A (u3_mem_b0_b_102 ), .B (n_3812), .S0 (n_8700), .Y(n_9388));
MX2X1 g34119(.A (u3_mem_b0_b_103 ), .B (n_3606), .S0 (n_8700), .Y(n_8724));
MX2X1 g34116(.A (u3_mem_b0_b ), .B (n_3808), .S0 (n_7423), .Y(n_8253));
MX2X1 g34117(.A (u3_mem_b0_b_100 ), .B (n_3809), .S0 (n_8700), .Y(n_8725));
MX2X1 g34114(.A (u7_mem_b0_b_98 ), .B (n_3625), .S0 (n_7493), .Y(n_8726));
MX2X1 g34115(.A (u7_mem_b0_b_99 ), .B (n_3626), .S0 (n_7493), .Y(n_9389));
MX2X1 g34112(.A (u7_mem_b0_b_96 ), .B (n_3631), .S0 (n_7493), .Y(n_8727));
MX2X1 g34113(.A (u7_mem_b0_b_97 ), .B (n_3623), .S0 (n_7493), .Y(n_9391));
MX2X1 g34110(.A (u7_mem_b0_b_94 ), .B (n_3619), .S0 (n_7493), .Y(n_9392));
MX2X1 g34111(.A (u7_mem_b0_b_95 ), .B (n_3620), .S0 (n_7493), .Y(n_8728));
NAND2X1 g36947(.A (n_1757), .B (n_1623), .Y (n_4017));
NAND2X1 g36946(.A (n_2528), .B (n_1235), .Y (n_4810));
NAND2X1 g34263(.A (u3_mem_b2_b_40 ), .B (n_8101), .Y (n_8138));
NAND2X1 g36945(.A (n_1629), .B (n_1625), .Y (n_4018));
NAND2X1 g36944(.A (n_1635), .B (n_1631), .Y (n_4019));
OAI21X1 g33588(.A0 (n_5085), .A1 (n_9336), .B0 (n_7965), .Y (n_9337));
OAI21X1 g33589(.A0 (n_5084), .A1 (n_9333), .B0 (n_7964), .Y (n_9335));
OAI21X1 g33858(.A0 (n_4311), .A1 (n_8981), .B0 (n_7667), .Y (n_8999));
OAI21X1 g33859(.A0 (n_4529), .A1 (n_8948), .B0 (n_7666), .Y (n_8998));
XOR2X1 g35491(.A (u2_res_cnt_b3_b ), .B (n_1278), .Y (n_4101));
OAI21X1 g33852(.A0 (n_4501), .A1 (n_9038), .B0 (n_7673), .Y (n_9005));
OAI21X1 g33853(.A0 (n_4510), .A1 (n_9036), .B0 (n_7672), .Y (n_9004));
OAI21X1 g33850(.A0 (n_4313), .A1 (n_9036), .B0 (n_7674), .Y (n_9008));
OAI21X1 g33851(.A0 (n_4496), .A1 (n_9043), .B0 (n_8078), .Y (n_9007));
OAI21X1 g33856(.A0 (n_4481), .A1 (n_9010), .B0 (n_7669), .Y (n_9001));
OAI21X1 g33857(.A0 (n_4312), .A1 (n_9010), .B0 (n_7668), .Y (n_9000));
OAI21X1 g33854(.A0 (n_4506), .A1 (n_9055), .B0 (n_7671), .Y (n_9003));
OAI21X1 g33855(.A0 (n_4516), .A1 (n_9034), .B0 (n_7670), .Y (n_9002));
NOR2X1 g39302(.A (n_5102), .B (n_2729), .Y (n_3295));
MX2X1 g35493(.A (u26_cnt_b1_b ), .B (n_794), .S0 (n_5624), .Y(n_5626));
MX2X1 g35494(.A (u26_cnt_b2_b ), .B (n_1821), .S0 (n_5624), .Y(n_5625));
AOI21X1 g38241(.A0 (u3_mem_b2_b_31 ), .A1 (n_4533), .B0 (n_2131), .Y(n_4394));
NAND2X1 g31727(.A (n_5498), .B (n_10385), .Y (n_10348));
NAND2X1 g36962(.A (n_1582), .B (n_1602), .Y (n_4007));
AOI21X1 g35497(.A0 (i3_re), .A1 (u9_rp_b0_b ), .B0 (n_6714), .Y(n_7143));
NAND2X1 g31724(.A (n_5492), .B (n_10376), .Y (n_10351));
NAND2X1 g39303(.A (n_2325), .B (in_slt_441), .Y (n_2326));
NAND2X1 g34644(.A (u6_mem_b2_b_29 ), .B (n_7758), .Y (n_7781));
NAND2X1 g31725(.A (n_5500), .B (n_10376), .Y (n_10350));
NAND2X1 g31722(.A (n_162), .B (n_10010), .Y (n_9975));
OAI21X1 g31051(.A0 (n_5293), .A1 (n_10450), .B0 (n_9986), .Y(n_10674));
INVX8 g40754(.A (n_1432), .Y (n_3316));
NAND2X1 g31720(.A (n_5488), .B (n_10385), .Y (n_10354));
NAND2X1 g31721(.A (n_5490), .B (n_10391), .Y (n_10353));
OAI21X1 g32989(.A0 (n_7327), .A1 (n_7175), .B0 (n_9885), .Y(n_12018));
OAI21X1 g32988(.A0 (n_7277), .A1 (n_7199), .B0 (n_9885), .Y(n_11676));
NAND2X1 g32987(.A (n_8175), .B (n_8673), .Y (n_9455));
AOI21X1 g32986(.A0 (n_7440), .A1 (n_7441), .B0 (n_8205), .Y (n_8206));
AOI21X1 g32985(.A0 (n_7381), .A1 (n_7382), .B0 (n_7524), .Y (n_7525));
AOI21X1 g32984(.A0 (n_7384), .A1 (n_7385), .B0 (n_7526), .Y (n_7527));
NAND2X1 g32983(.A (n_8177), .B (n_8674), .Y (n_9456));
NAND2X1 g32982(.A (n_8181), .B (n_8675), .Y (n_9457));
NAND2X1 g32981(.A (n_8178), .B (n_8676), .Y (n_9458));
NAND2X1 g32980(.A (n_8179), .B (n_8677), .Y (n_9459));
NAND2X1 g34642(.A (u6_mem_b2_b_46 ), .B (n_7758), .Y (n_7783));
INVX1 g39503(.A (n_4743), .Y (n_3137));
NOR2X1 g37139(.A (n_2599), .B (n_1263), .Y (n_2600));
MX2X1 g38618(.A (u4_mem_b0_b_108 ), .B (wb_din_678), .S0 (n_3765), .Y(n_3784));
NAND2X1 g32679(.A (n_335), .B (n_10645), .Y (n_11957));
AOI21X1 g32678(.A0 (n_6227), .A1 (n_6225), .B0 (n_9876), .Y(n_10633));
AOI21X1 g40386(.A0 (u4_rp_b3_b ), .A1 (u4_wp_b2_b ), .B0 (n_441), .Y(n_1001));
XOR2X1 g40387(.A (n_886), .B (n_657), .Y (n_2645));
XOR2X1 g40380(.A (n_614), .B (n_868), .Y (n_2646));
AOI22X1 g40381(.A0 (n_496), .A1 (n_1255), .B0 (u6_rp_b3_b ), .B1(u6_wp_b2_b ), .Y (n_1256));
AOI22X1 g40383(.A0 (n_457), .A1 (n_1443), .B0 (u7_rp_b3_b ), .B1(u7_wp_b2_b ), .Y (n_1444));
NAND2X1 g32671(.A (n_134), .B (n_10645), .Y (n_11955));
NAND2X1 g32670(.A (n_186), .B (n_10645), .Y (n_11979));
NAND2X1 g32673(.A (n_163), .B (n_10645), .Y (n_11975));
NAND2X1 g32672(.A (n_254), .B (n_10645), .Y (n_11991));
NAND2X1 g32675(.A (n_399), .B (n_10645), .Y (n_10636));
NAND2X1 g32674(.A (n_230), .B (n_10605), .Y (n_11734));
AOI21X1 g32677(.A0 (n_6784), .A1 (n_5845), .B0 (n_9876), .Y(n_10634));
NAND2X1 g32676(.A (n_299), .B (n_10645), .Y (n_11973));
NAND4X1 g37000(.A (n_12819), .B (n_1415), .C (n_12820), .D (n_2416),.Y (n_6224));
INVX1 g37003(.A (n_5841), .Y (n_5548));
NAND4X1 g37002(.A (n_12821), .B (n_2855), .C (n_12822), .D (n_2376),.Y (n_6226));
INVX1 g37005(.A (n_5837), .Y (n_5547));
NAND4X1 g37004(.A (n_11709), .B (n_11710), .C (n_2276), .D (n_2413),.Y (n_5841));
MX2X1 g38767(.A (u7_mem_b0_b_111 ), .B (wb_din_681), .S0 (n_3622), .Y(n_3568));
NAND4X1 g37006(.A (n_11711), .B (n_11712), .C (n_2272), .D (n_2398),.Y (n_5837));
NAND4X1 g37009(.A (n_11660), .B (n_11661), .C (n_2355), .D (n_3529),.Y (n_6248));
INVX1 g37008(.A (n_6248), .Y (n_5701));
AOI21X1 g38345(.A0 (u5_mem_b3_b_138 ), .A1 (n_4996), .B0 (n_3133), .Y(n_4992));
AOI21X1 g38344(.A0 (u5_mem_b3_b_137 ), .A1 (n_5000), .B0 (n_3154), .Y(n_4993));
AND2X1 g36608(.A (n_5384), .B (n_1779), .Y (n_5797));
NAND2X1 g36609(.A (n_6144), .B (n_634), .Y (n_6145));
NAND2X1 g36358(.A (n_6783), .B (n_6821), .Y (n_6820));
NAND2X1 g36359(.A (n_6226), .B (n_6821), .Y (n_6305));
NAND2X1 g36604(.A (n_6147), .B (n_6118), .Y (n_12047));
NAND2X1 g36357(.A (n_6224), .B (n_6821), .Y (n_6307));
NAND2X1 g36606(.A (n_12514), .B (n_6773), .Y (n_6146));
INVX4 g36607(.A (n_5797), .Y (n_7353));
NAND2X1 g36600(.A (n_6153), .B (n_6152), .Y (n_6154));
NAND2X1 g36602(.A (n_6150), .B (n_12664), .Y (n_6151));
NAND2X1 g36351(.A (n_6786), .B (n_6821), .Y (n_6822));
AOI22X1 g37318(.A0 (n_4729), .A1 (n_8199), .B0 (n_5591), .B1(n_4736), .Y (n_4737));
AOI21X1 g38341(.A0 (u5_mem_b3_b_134 ), .A1 (n_4996), .B0 (n_2932), .Y(n_4997));
NAND2X1 g39089(.A (u8_mem_b1_b_69 ), .B (n_12295), .Y (n_11452));
AOI21X1 g38340(.A0 (u5_mem_b3_b_133 ), .A1 (n_5000), .B0 (n_2739), .Y(n_4998));
AOI22X1 g37747(.A0 (n_215), .A1 (n_2530), .B0 (n_2545), .B1 (n_2544),.Y (n_2547));
NOR2X1 g40143(.A (n_2801), .B (n_2137), .Y (n_2092));
NAND2X1 g39309(.A (u7_mem_b1_b_89 ), .B (n_4130), .Y (n_4203));
MX2X1 g38589(.A (u8_mem_b0_b_109 ), .B (wb_din_679), .S0 (n_3826), .Y(n_3827));
MX2X1 g38588(.A (u8_mem_b0_b_91 ), .B (wb_din_661), .S0 (n_3826), .Y(n_3828));
MX2X1 g38585(.A (u8_mem_b0_b_93 ), .B (wb_din_663), .S0 (n_3826), .Y(n_3832));
MX2X1 g38584(.A (u8_mem_b0_b_112 ), .B (wb_din_682), .S0 (n_3826), .Y(n_3833));
MX2X1 g38587(.A (u8_mem_b0_b_110 ), .B (wb_din_680), .S0 (n_3826), .Y(n_3830));
MX2X1 g38586(.A (u8_mem_b0_b_111 ), .B (wb_din_681), .S0 (n_3826), .Y(n_3831));
MX2X1 g38581(.A (u8_mem_b0_b_94 ), .B (wb_din_664), .S0 (n_3826), .Y(n_3837));
MX2X1 g38580(.A (u8_mem_b0_b_114 ), .B (wb_din_684), .S0 (n_3826), .Y(n_3838));
MX2X1 g38583(.A (u3_mem_b0_b_112 ), .B (wb_din_682), .S0 (n_858), .Y(n_3834));
MX2X1 g38582(.A (u8_mem_b0_b_113 ), .B (wb_din_683), .S0 (n_3826), .Y(n_3836));
NOR2X1 g40145(.A (n_2749), .B (n_2748), .Y (n_2750));
OAI21X1 g33733(.A0 (n_5113), .A1 (n_9182), .B0 (n_7796), .Y (n_9152));
NOR2X1 g40148(.A (n_2773), .B (n_2741), .Y (n_2747));
NOR2X1 g40218(.A (n_2081), .B (n_2735), .Y (n_2030));
AOI21X1 g30834(.A0 (n_11990), .A1 (n_11991), .B0 (n_11086), .Y(n_11087));
INVX2 g41381(.A (n_12678), .Y (n_1397));
INVX4 g41380(.A (n_1397), .Y (n_3259));
INVX8 g41384(.A (n_1396), .Y (n_6594));
NAND2X1 g39505(.A (n_11798), .B (u8_mem_b0_b_116 ), .Y (n_3136));
INVX1 g41389(.A (n_1067), .Y (n_1396));
MX2X1 g31379(.A (u11_din_tmp_43), .B (in_slt_446), .S0 (n_10103), .Y(n_10104));
MX2X1 g31378(.A (u11_din_tmp_42), .B (in_slt_445), .S0 (n_10103), .Y(n_10105));
MX2X1 g31375(.A (u11_din_tmp_54), .B (in_slt_457), .S0 (n_10103), .Y(n_10110));
MX2X1 g31374(.A (u11_din_tmp_53), .B (in_slt_456), .S0 (n_10103), .Y(n_10111));
MX2X1 g31377(.A (u11_din_tmp_56), .B (in_slt_459), .S0 (n_10103), .Y(n_10106));
MX2X1 g31376(.A (u11_din_tmp_55), .B (in_slt_458), .S0 (n_10103), .Y(n_10108));
MX2X1 g31371(.A (u11_din_tmp1), .B (in_slt_444), .S0 (n_10103), .Y(n_10115));
MX2X1 g31370(.A (u10_din_tmp_50), .B (in_slt_431), .S0 (n_9860), .Y(n_9862));
MX2X1 g31373(.A (u11_din_tmp_52), .B (in_slt_455), .S0 (n_10103), .Y(n_10112));
MX2X1 g31372(.A (u11_din_tmp_51), .B (in_slt_454), .S0 (n_10103), .Y(n_10114));
AOI21X1 g38025(.A0 (u3_mem_b2_b_29 ), .A1 (n_4533), .B0 (n_1963), .Y(n_4526));
AOI22X1 g37919(.A0 (u11_din_tmp_49), .A1 (n_4560), .B0 (n_4097), .B1(in_slt_450), .Y (n_4561));
AOI22X1 g37917(.A0 (u11_din_tmp_48), .A1 (n_4560), .B0 (n_4097), .B1(in_slt_449), .Y (n_4563));
NAND2X1 g37916(.A (n_4200), .B (n_3225), .Y (n_5463));
AOI22X1 g37915(.A0 (n_6656), .A1 (n_1859), .B0 (n_6620), .B1(n_1760), .Y (n_1848));
AOI22X1 g37913(.A0 (u11_din_tmp_47), .A1 (n_4560), .B0 (n_4097), .B1(in_slt_448), .Y (n_4565));
AOI22X1 g37911(.A0 (u11_din_tmp_46), .A1 (n_4560), .B0 (n_4097), .B1(in_slt_447), .Y (n_4566));
AOI22X1 g37910(.A0 (u11_din_tmp_45), .A1 (n_4560), .B0 (n_4097), .B1(in_slt_446), .Y (n_4567));
MX2X1 g33209(.A (u13_intm_r_b27_b ), .B (wb_din_687), .S0 (n_8519), .Y(n_8498));
MX2X1 g33208(.A (u13_intm_r_b26_b ), .B (wb_din_686), .S0 (n_8519), .Y(n_8500));
MX2X1 g33207(.A (u13_intm_r_b25_b ), .B (wb_din_685), .S0 (n_8519), .Y(n_8502));
MX2X1 g33206(.A (u13_intm_r_b24_b ), .B (wb_din_684), .S0 (n_8519), .Y(n_8504));
MX2X1 g33205(.A (u13_intm_r_b23_b ), .B (wb_din_683), .S0 (n_8519), .Y(n_8505));
MX2X1 g33204(.A (u13_intm_r_b22_b ), .B (wb_din_682), .S0 (n_8519), .Y(n_8506));
MX2X1 g33203(.A (u13_intm_r_b21_b ), .B (wb_din_681), .S0 (n_8519), .Y(n_8507));
MX2X1 g33202(.A (u13_intm_r_b20_b ), .B (wb_din_680), .S0 (n_8519), .Y(n_8508));
MX2X1 g33201(.A (u13_intm_r_b1_b ), .B (wb_din_661), .S0 (n_8519), .Y(n_8509));
MX2X1 g33200(.A (u13_intm_r_b19_b ), .B (wb_din_679), .S0 (n_8519), .Y(n_8510));
INVX1 g42128(.A (u9_mem_b1_b_119 ), .Y (n_6949));
INVX1 g42129(.A (u9_mem_b3_b_83 ), .Y (n_5367));
INVX1 g42122(.A (u10_mem_b3_b_63 ), .Y (n_6562));
INVX1 g42120(.A (u9_mem_b2_b_115 ), .Y (n_345));
INVX1 g42124(.A (u11_mem_b0_b ), .Y (n_6377));
INVX1 g42125(.A (u9_mem_b3_b_67 ), .Y (n_6617));
MX2X1 g35982(.A (n_6956), .B (n_6925), .S0 (n_5730), .Y (n_6957));
MX2X1 g35983(.A (n_6656), .B (n_6646), .S0 (n_4783), .Y (n_6657));
MX2X1 g35980(.A (n_5987), .B (n_6026), .S0 (n_6649), .Y (n_6027));
MX2X1 g35981(.A (n_6486), .B (n_6658), .S0 (n_6649), .Y (n_6659));
MX2X1 g35986(.A (n_5993), .B (n_6023), .S0 (n_6649), .Y (n_6024));
MX2X1 g35987(.A (n_6952), .B (n_6951), .S0 (n_6908), .Y (n_6953));
MX2X1 g35984(.A (n_6654), .B (n_6637), .S0 (n_4783), .Y (n_6655));
MX2X1 g35985(.A (n_6954), .B (n_6952), .S0 (n_4783), .Y (n_6955));
NOR2X1 g39959(.A (n_2829), .B (n_1488), .Y (n_1556));
MX2X1 g35988(.A (n_6949), .B (n_6920), .S0 (n_969), .Y (n_6950));
MX2X1 g35989(.A (n_6947), .B (n_6891), .S0 (n_4783), .Y (n_6948));
NOR2X1 g40048(.A (n_2836), .B (n_2804), .Y (n_2805));
NOR2X1 g39305(.A (n_3486), .B (n_2831), .Y (n_3292));
AOI21X1 g31656(.A0 (n_7288), .A1 (n_1208), .B0 (n_9503), .Y (n_9504));
BUFX3 g35188(.A (o8_we), .Y (n_7402));
INVX1 g35181(.A (n_7402), .Y (n_9038));
INVX2 g35187(.A (n_7402), .Y (n_9034));
INVX1 g35185(.A (n_7402), .Y (n_9010));
NAND2X1 g34857(.A (u8_mem_b2_b_43 ), .B (n_7976), .Y (n_7577));
NAND2X1 g34856(.A (u3_mem_b1_b_78 ), .B (n_8141), .Y (n_7578));
NAND2X1 g34855(.A (u8_mem_b2_b_42 ), .B (n_7976), .Y (n_7579));
NAND2X1 g34854(.A (u8_mem_b2_b_47 ), .B (n_7976), .Y (n_7580));
NAND2X1 g34852(.A (u8_mem_b2_b_40 ), .B (n_7976), .Y (n_7582));
NAND2X1 g34851(.A (u8_mem_b2_b_38 ), .B (n_7976), .Y (n_7583));
NAND2X1 g34850(.A (u8_mem_b2_b ), .B (n_7976), .Y (n_7584));
NAND2X1 g34859(.A (u3_mem_b1_b_60 ), .B (n_8101), .Y (n_7575));
NAND2X1 g34858(.A (u8_mem_b2_b_44 ), .B (n_7976), .Y (n_7576));
AOI21X1 g30135(.A0 (n_5964), .A1 (n_11131), .B0 (n_11006), .Y(n_11518));
AOI21X1 g30137(.A0 (n_5636), .A1 (n_11126), .B0 (n_11004), .Y(n_11516));
NAND2X1 g35450(.A (n_7298), .B (n_6743), .Y (n_7451));
MX2X1 g30138(.A (n_4801), .B (n_10095), .S0 (n_10992), .Y (n_10969));
MX2X1 g30139(.A (n_2594), .B (n_10094), .S0 (n_10985), .Y (n_10968));
NAND2X1 g35328(.A (n_6720), .B (n_11600), .Y (n_7380));
NAND2X1 g35329(.A (n_7030), .B (n_11772), .Y (n_7439));
NAND4X1 g36982(.A (n_11707), .B (n_11708), .C (n_2282), .D (n_2447),.Y (n_5853));
INVX1 g36981(.A (n_5853), .Y (n_5552));
NAND4X1 g36980(.A (n_3091), .B (n_2925), .C (n_4246), .D (n_1861), .Y(n_6779));
INVX1 g36987(.A (n_5851), .Y (n_5551));
NAND2X1 g36986(.A (n_1570), .B (n_1689), .Y (n_4003));
NAND4X1 g36985(.A (n_3078), .B (n_2868), .C (n_2287), .D (n_2433), .Y(n_5805));
NAND4X1 g36984(.A (n_11697), .B (n_11698), .C (n_4164), .D (n_2452),.Y (n_6786));
NAND4X1 g36988(.A (n_11699), .B (n_11700), .C (n_2278), .D (n_2424),.Y (n_5851));
NAND2X1 g34581(.A (u5_mem_b3_b_125 ), .B (n_7870), .Y (n_7845));
NAND2X1 g34580(.A (u5_mem_b3_b_124 ), .B (n_7870), .Y (n_7846));
NAND2X1 g34583(.A (u5_mem_b3_b_127 ), .B (n_7870), .Y (n_7843));
NAND2X1 g34582(.A (u5_mem_b3_b_126 ), .B (n_7870), .Y (n_7844));
NAND2X1 g34585(.A (u5_mem_b3_b_129 ), .B (n_7870), .Y (n_7841));
NAND2X1 g34584(.A (u5_mem_b3_b_128 ), .B (n_7870), .Y (n_7842));
NAND2X1 g34587(.A (u8_mem_b1_b_75 ), .B (n_7976), .Y (n_7839));
NAND2X1 g34586(.A (u5_mem_b3_b_130 ), .B (n_7870), .Y (n_7840));
NOR2X1 g34589(.A (n_798), .B (n_7870), .Y (n_8224));
NAND2X1 g34588(.A (u8_mem_b3_b_131 ), .B (n_7976), .Y (n_7838));
INVX8 g32866(.A (n_9726), .Y (n_10315));
INVX4 g32867(.A (n_9676), .Y (n_9726));
NAND2X1 g36496(.A (n_6816), .B (n_5853), .Y (n_5854));
MX2X1 g34003(.A (u4_mem_b0_b_92 ), .B (n_3761), .S0 (n_7499), .Y(n_8817));
NAND2X1 g36493(.A (n_3561), .B (n_1291), .Y (n_4835));
OR2X1 g19(.A (n_1374), .B (n_12340), .Y (n_11841));
OR2X1 g18(.A (n_12687), .B (n_12534), .Y (n_12339));
OAI21X1 g16(.A0 (n_11904), .A1 (n_11504), .B0 (n_11905), .Y(n_11906));
INVX2 g12(.A (u7_rp_b1_b ), .Y (n_12330));
INVX2 g11(.A (n_12330), .Y (n_12331));
INVX2 g10(.A (u7_rp_b2_b ), .Y (n_12332));
NOR2X1 g39069(.A (n_3089), .B (n_2755), .Y (n_3478));
OAI21X1 g33445(.A0 (n_4528), .A1 (n_8911), .B0 (n_8131), .Y (n_8418));
OAI21X1 g33444(.A0 (n_3861), .A1 (n_8457), .B0 (n_7833), .Y (n_8419));
OAI21X1 g33447(.A0 (n_4296), .A1 (n_8097), .B0 (n_7723), .Y (n_8415));
OAI21X1 g33446(.A0 (n_3877), .A1 (n_8449), .B0 (n_7836), .Y (n_8416));
NAND2X1 g34321(.A (u8_mem_b2_b_45 ), .B (n_7976), .Y (n_8076));
NAND2X1 g34320(.A (u3_mem_b3_b_124 ), .B (n_8101), .Y (n_8077));
NAND2X1 g34323(.A (u3_mem_b3_b_128 ), .B (n_8141), .Y (n_8074));
OAI21X1 g33442(.A0 (n_4325), .A1 (n_8856), .B0 (n_8136), .Y (n_8421));
OAI21X1 g33449(.A0 (n_4486), .A1 (n_8856), .B0 (n_8129), .Y (n_8412));
OAI21X1 g33448(.A0 (n_4277), .A1 (n_8898), .B0 (n_8126), .Y (n_8413));
NAND2X1 g36319(.A (n_6807), .B (n_6824), .Y (n_11539));
OAI21X1 g45800(.A0 (n_12520), .A1 (n_12521), .B0 (n_12609), .Y(n_12813));
MX2X1 g37214(.A (u10_mem_b2_b_111 ), .B (n_5287), .S0 (n_5341), .Y(n_5378));
NAND2X1 g34732(.A (u7_mem_b1_b_83 ), .B (n_7651), .Y (n_7702));
AOI21X1 g37216(.A0 (n_5522), .A1 (n_6649), .B0 (n_4635), .Y (n_5523));
MX2X1 g37217(.A (u10_mem_b1_b_146 ), .B (n_4751), .S0 (n_6475), .Y(n_4792));
AOI21X1 g37210(.A0 (n_5524), .A1 (n_6649), .B0 (n_4636), .Y (n_5525));
MX2X1 g37211(.A (u10_mem_b2_b_107 ), .B (n_5292), .S0 (n_5341), .Y(n_5380));
MX2X1 g37212(.A (u10_mem_b2_b_108 ), .B (n_4745), .S0 (n_5424), .Y(n_4793));
NAND2X1 g34733(.A (u7_mem_b1_b_84 ), .B (n_7651), .Y (n_7701));
NAND2X1 g37748(.A (n_3555), .B (n_3493), .Y (n_4595));
NAND2X1 g37749(.A (n_2443), .B (n_2316), .Y (n_3914));
MX2X1 g37218(.A (u9_mem_b1_b_138 ), .B (n_4778), .S0 (n_5730), .Y(n_4791));
NAND2X1 g34730(.A (u7_mem_b1_b_81 ), .B (n_7651), .Y (n_7704));
XOR2X1 g38248(.A (n_1255), .B (n_5059), .Y (n_4389));
AOI21X1 g38249(.A0 (u6_mem_b3_b_130 ), .A1 (n_5100), .B0 (n_2777), .Y(n_5058));
OAI21X1 g33052(.A0 (n_7328), .A1 (n_7202), .B0 (n_9885), .Y(n_11988));
OAI21X1 g33053(.A0 (n_7230), .A1 (n_7079), .B0 (n_12161), .Y(n_12793));
OAI21X1 g33050(.A0 (n_7203), .A1 (n_7081), .B0 (n_12161), .Y(n_12064));
OAI21X1 g33057(.A0 (n_7227), .A1 (n_7076), .B0 (n_10481), .Y(n_11749));
OAI21X1 g33054(.A0 (n_7306), .A1 (n_6987), .B0 (n_12161), .Y(n_10188));
OAI21X1 g33055(.A0 (n_7271), .A1 (n_7095), .B0 (n_10481), .Y(n_11743));
INVX1 g34880(.A (n_9710), .Y (n_9689));
OAI21X1 g33059(.A0 (n_7225), .A1 (n_7073), .B0 (n_12689), .Y(n_10504));
NOR2X1 g34882(.A (n_7285), .B (n_2595), .Y (n_7438));
NAND2X1 g34883(.A (n_9470), .B (n_9579), .Y (n_9580));
NAND2X1 g34369(.A (u4_mem_b1_b_84 ), .B (n_7984), .Y (n_8033));
NAND2X1 g34739(.A (u7_mem_b1_b_88 ), .B (n_7651), .Y (n_7695));
NOR2X1 g40235(.A (n_938), .B (n_2686), .Y (n_2019));
NAND2X1 g39228(.A (u3_mem_b1_b_81 ), .B (n_3316), .Y (n_3354));
NOR2X1 g39588(.A (n_3453), .B (n_2716), .Y (n_3079));
OAI21X1 g33401(.A0 (n_4489), .A1 (n_8464), .B0 (n_8173), .Y (n_8475));
AOI22X1 g33400(.A0 (n_4299), .A1 (n_7493), .B0 (n_7651), .B1(u7_wp_b2_b ), .Y (n_8476));
OAI21X1 g33403(.A0 (n_4490), .A1 (n_8894), .B0 (n_8070), .Y (n_8473));
NOR2X1 g41596(.A (n_751), .B (n_706), .Y (n_707));
INVX4 g41594(.A (n_5059), .Y (n_1509));
OAI21X1 g33405(.A0 (n_5158), .A1 (n_8911), .B0 (n_8169), .Y (n_8471));
OR2X1 g41598(.A (n_1372), .B (n_2485), .Y (n_1373));
NAND2X1 g34364(.A (u4_mem_b1_b_80 ), .B (n_7984), .Y (n_8037));
MX2X1 g36165(.A (n_5957), .B (n_6014), .S0 (n_6341), .Y (n_5958));
AOI21X1 g30897(.A0 (n_11635), .A1 (n_11636), .B0 (n_11036), .Y(n_11021));
MX2X1 g36167(.A (n_6360), .B (n_6459), .S0 (n_6359), .Y (n_6361));
MX2X1 g36166(.A (n_6363), .B (n_6465), .S0 (n_6359), .Y (n_6364));
MX2X1 g36161(.A (n_6372), .B (n_6478), .S0 (n_6359), .Y (n_6373));
OAI21X1 g33407(.A0 (n_4530), .A1 (n_8464), .B0 (n_8168), .Y (n_8469));
MX2X1 g36163(.A (n_6368), .B (n_6514), .S0 (n_6359), .Y (n_6369));
AOI21X1 g35604(.A0 (n_6271), .A1 (n_5764), .B0 (n_7267), .Y (n_7258));
NAND2X1 g34366(.A (u4_mem_b1_b_82 ), .B (n_7984), .Y (n_8035));
MX2X1 g36169(.A (n_5953), .B (n_5993), .S0 (n_6359), .Y (n_5954));
AOI21X1 g35607(.A0 (n_5924), .A1 (n_6113), .B0 (n_7256), .Y (n_7254));
AOI21X1 g35606(.A0 (n_5925), .A1 (n_6114), .B0 (n_7256), .Y (n_7255));
INVX1 g42719(.A (n_459), .Y (n_862));
NAND2X1 g39586(.A (in_slt_412), .B (n_3415), .Y (n_3081));
AOI21X1 g35600(.A0 (n_5888), .A1 (n_5931), .B0 (n_12604), .Y(n_7126));
INVX2 g40971(.A (n_930), .Y (n_1158));
AOI21X1 g31748(.A0 (n_9536), .A1 (n_10518), .B0 (n_676), .Y(n_10798));
AOI21X1 g31749(.A0 (n_2360), .A1 (n_4834), .B0 (n_11892), .Y(n_9969));
AOI21X1 g31744(.A0 (n_9541), .A1 (n_12149), .B0 (n_540), .Y (n_9972));
INVX1 g31745(.A (n_9970), .Y (n_10343));
AOI21X1 g31746(.A0 (n_9538), .A1 (n_12609), .B0 (n_665), .Y (n_9970));
INVX1 g31747(.A (n_10798), .Y (n_10906));
AOI22X1 g31740(.A0 (n_7520), .A1 (n_8207), .B0 (n_565), .B1 (n_7434),.Y (n_9446));
INVX1 g31741(.A (n_10799), .Y (n_10907));
AOI21X1 g31742(.A0 (n_9543), .A1 (n_12689), .B0 (n_616), .Y(n_10799));
NOR2X1 g35669(.A (n_5444), .B (n_1274), .Y (n_6061));
AOI21X1 g35668(.A0 (n_12046), .A1 (n_12047), .B0 (n_12640), .Y(n_7203));
NOR2X1 g30839(.A (n_10989), .B (n_11086), .Y (n_11148));
NOR2X1 g30838(.A (n_10991), .B (n_11086), .Y (n_11149));
AOI21X1 g35849(.A0 (n_2584), .A1 (n_5273), .B0 (n_7353), .Y (n_7109));
AOI21X1 g35848(.A0 (n_2585), .A1 (n_5274), .B0 (n_7353), .Y (n_7045));
AOI21X1 g30835(.A0 (n_11974), .A1 (n_11975), .B0 (n_11083), .Y(n_11085));
AOI21X1 g35662(.A0 (n_6278), .A1 (n_5767), .B0 (n_7214), .Y (n_7208));
AOI21X1 g30837(.A0 (n_11972), .A1 (n_11973), .B0 (n_5827), .Y(n_11082));
AOI21X1 g30836(.A0 (n_10636), .A1 (n_10523), .B0 (n_11083), .Y(n_11084));
AOI21X1 g30831(.A0 (n_11952), .A1 (n_11953), .B0 (n_11083), .Y(n_11092));
AOI21X1 g30830(.A0 (n_11968), .A1 (n_11969), .B0 (n_1870), .Y(n_11093));
AOI21X1 g30833(.A0 (n_11954), .A1 (n_11955), .B0 (n_5827), .Y(n_11089));
AOI21X1 g30832(.A0 (n_11978), .A1 (n_11979), .B0 (n_11083), .Y(n_11091));
NAND2X1 g38835(.A (u4_mem_b3_b_149 ), .B (n_3556), .Y (n_3548));
AOI22X1 g37822(.A0 (n_5966), .A1 (n_1839), .B0 (n_6002), .B1(n_1316), .Y (n_1612));
INVX1 g35542(.A (i4_full), .Y (n_631));
AOI22X1 g37821(.A0 (n_275), .A1 (n_1575), .B0 (n_5496), .B1 (n_1831),.Y (n_1613));
AOI22X1 g37356(.A0 (n_5272), .A1 (u13_intm_r_b8_b ), .B0 (n_5277), .B1(crac_din_699), .Y (n_5258));
NAND2X1 g45681(.A (dma_req_o_b7_b), .B (n_12375), .Y (n_12377));
NAND2X1 g38832(.A (u3_mem_b3_b_144 ), .B (n_2463), .Y (n_2446));
NAND2X1 g36512(.A (n_5844), .B (n_1297), .Y (n_5845));
OAI21X1 g35933(.A0 (n_5667), .A1 (n_7063), .B0 (n_5812), .Y (n_7065));
OAI21X1 g35932(.A0 (n_5677), .A1 (n_7077), .B0 (n_6263), .Y (n_7066));
NAND2X1 g38839(.A (u8_mem_b3_b_143 ), .B (n_2468), .Y (n_2445));
OAI21X1 g35931(.A0 (n_5534), .A1 (n_7063), .B0 (n_5814), .Y (n_6984));
NAND2X1 g38838(.A (u7_mem_b3_b_131 ), .B (n_1538), .Y (n_1545));
XOR2X1 g35492(.A (u2_to_cnt_b3_b ), .B (n_1276), .Y (n_4100));
OAI21X1 g35930(.A0 (n_5698), .A1 (n_7077), .B0 (n_6187), .Y (n_7067));
OAI21X1 g35937(.A0 (n_5530), .A1 (n_6981), .B0 (n_5810), .Y (n_6982));
OAI21X1 g35936(.A0 (n_5668), .A1 (n_7077), .B0 (n_6173), .Y (n_7062));
NAND2X1 g45668(.A (n_12622), .B (u6_mem_b3_b_137 ), .Y (n_12362));
OAI21X1 g35935(.A0 (n_5532), .A1 (n_6981), .B0 (n_5808), .Y (n_6983));
NAND2X1 g45669(.A (u6_mem_b1_b_75 ), .B (n_12169), .Y (n_12363));
OAI21X1 g35934(.A0 (n_5533), .A1 (n_7063), .B0 (n_6183), .Y (n_7064));
MX2X1 g34138(.A (u8_mem_b0_b_91 ), .B (n_3828), .S0 (n_7490), .Y(n_8708));
MX2X1 g34139(.A (u3_mem_b0_b_111 ), .B (n_3593), .S0 (n_8700), .Y(n_9380));
INVX1 g39907(.A (n_5292), .Y (n_4111));
MX2X1 g34130(.A (u8_mem_b0_b_104 ), .B (n_3600), .S0 (n_7490), .Y(n_8717));
MX2X1 g34131(.A (u8_mem_b0_b_105 ), .B (n_3824), .S0 (n_7490), .Y(n_8715));
MX2X1 g34132(.A (u8_mem_b0_b_106 ), .B (n_3599), .S0 (n_7490), .Y(n_8714));
MX2X1 g34133(.A (u3_mem_b0_b_91 ), .B (n_3598), .S0 (n_8700), .Y(n_9382));
MX2X1 g34134(.A (u8_mem_b0_b_107 ), .B (n_3825), .S0 (n_7490), .Y(n_9381));
MX2X1 g34135(.A (u8_mem_b0_b_108 ), .B (n_3596), .S0 (n_7490), .Y(n_8713));
MX2X1 g34136(.A (u3_mem_b0_b_110 ), .B (n_3595), .S0 (n_8700), .Y(n_8711));
MX2X1 g34137(.A (u8_mem_b0_b_109 ), .B (n_3827), .S0 (n_7490), .Y(n_8709));
NOR2X1 g40357(.A (n_2025), .B (n_2712), .Y (n_1942));
NAND2X1 g39905(.A (n_12679), .B (u5_mem_b0_b_112 ), .Y (n_2889));
INVX1 g41547(.A (n_2419), .Y (n_1377));
NOR2X1 g40356(.A (n_1226), .B (n_2763), .Y (n_2656));
NAND3X1 g39270(.A (u3_mem_b0_b_91 ), .B (n_814), .C (n_1924), .Y(n_1487));
NOR2X1 g39271(.A (u10_mem_b1_b_138 ), .B (n_2364), .Y (n_2335));
NAND2X1 g39744(.A (n_12825), .B (u3_mem_b0_b_120 ), .Y (n_2984));
NAND2X1 g39745(.A (u4_mem_b2_b_55 ), .B (n_12087), .Y (n_2983));
NAND2X1 g39746(.A (n_12679), .B (u5_mem_b0_b_118 ), .Y (n_2982));
NAND2X1 g39747(.A (u3_mem_b2_b_51 ), .B (n_3330), .Y (n_2981));
OR2X1 g39740(.A (n_1052), .B (u3_rp_b3_b ), .Y (n_2986));
NOR2X1 g39741(.A (n_3117), .B (n_2729), .Y (n_3053));
NOR2X1 g39742(.A (n_5138), .B (n_2681), .Y (n_2985));
NAND2X1 g39743(.A (u6_mem_b1_b_60 ), .B (n_12169), .Y (n_12820));
NOR2X1 g39273(.A (n_5138), .B (n_2772), .Y (n_3329));
NAND2X1 g39748(.A (n_12389), .B (u4_mem_b0_b_101 ), .Y (n_11654));
NAND2X1 g39749(.A (u4_mem_b1_b_90 ), .B (n_12270), .Y (n_4136));
NOR2X1 g40352(.A (n_2043), .B (n_2818), .Y (n_1944));
OAI21X1 g33875(.A0 (n_4887), .A1 (n_8981), .B0 (n_7649), .Y (n_8979));
OAI21X1 g33876(.A0 (n_4874), .A1 (n_8976), .B0 (n_7648), .Y (n_8978));
OAI21X1 g33877(.A0 (n_4886), .A1 (n_8976), .B0 (n_7647), .Y (n_8977));
OAI21X1 g33872(.A0 (n_4875), .A1 (n_8981), .B0 (n_7653), .Y (n_8983));
OAI21X1 g33873(.A0 (n_4888), .A1 (n_8981), .B0 (n_7652), .Y (n_8982));
INVX1 g42944(.A (n_8190), .Y (n_921));
OAI21X1 g33878(.A0 (n_4949), .A1 (n_8976), .B0 (n_7646), .Y (n_8975));
OAI21X1 g33879(.A0 (n_4962), .A1 (n_8976), .B0 (n_7645), .Y (n_8974));
AND2X1 g39057(.A (n_1225), .B (wb_addr_i_b4_b), .Y (n_3985));
AOI22X1 g37642(.A0 (n_345), .A1 (n_1835), .B0 (n_5347), .B1 (n_1760),.Y (n_1722));
NOR2X1 g39050(.A (n_3486), .B (n_2818), .Y (n_3487));
NAND2X1 g45667(.A (n_3474), .B (u6_mem_b2_b_44 ), .Y (n_12361));
NAND2X1 g39051(.A (u4_mem_b1_b_81 ), .B (n_12270), .Y (n_4236));
INVX1 g41844(.A (u10_mem_b3_b_80 ), .Y (n_5514));
AOI22X1 g37641(.A0 (n_2502), .A1 (n_1724), .B0 (n_1723), .B1(n_1859), .Y (n_1725));
INVX1 g41845(.A (u9_mem_b2_b_112 ), .Y (n_1700));
NOR2X1 g40358(.A (n_1016), .B (n_2864), .Y (n_2655));
AOI22X1 g37640(.A0 (n_346), .A1 (n_1835), .B0 (n_5367), .B1 (n_1760),.Y (n_1726));
AOI21X1 g38061(.A0 (u3_mem_b3_b_147 ), .A1 (n_5133), .B0 (n_3465), .Y(n_5129));
AOI21X1 g38067(.A0 (u8_mem_b2_b_44 ), .A1 (n_4499), .B0 (n_2153), .Y(n_4497));
AOI22X1 g37647(.A0 (n_2502), .A1 (n_6857), .B0 (n_6947), .B1(n_1859), .Y (n_1714));
AOI22X1 g37891(.A0 (n_3911), .A1 (in_slt_436), .B0 (n_2344), .B1(in_slt_434), .Y (n_2520));
MX2X1 g36015(.A (n_6612), .B (n_6566), .S0 (n_5341), .Y (n_6613));
AOI22X1 g37646(.A0 (n_2502), .A1 (n_1716), .B0 (n_1715), .B1(n_1859), .Y (n_1717));
NAND2X1 g32653(.A (n_113), .B (n_9931), .Y (n_9926));
NAND2X1 g32652(.A (n_101), .B (n_9931), .Y (n_9927));
NAND2X1 g32651(.A (n_261), .B (n_9931), .Y (n_9928));
NAND2X1 g32650(.A (n_300), .B (n_9931), .Y (n_9929));
AOI21X1 g32657(.A0 (n_5870), .A1 (n_5868), .B0 (n_9931), .Y (n_9921));
NAND2X1 g32656(.A (n_102), .B (n_9931), .Y (n_9922));
NAND2X1 g32655(.A (n_117), .B (n_9931), .Y (n_12836));
NAND2X1 g32654(.A (n_114), .B (n_9931), .Y (n_9925));
NAND2X1 g32659(.A (n_304), .B (n_9931), .Y (n_11999));
AOI21X1 g32658(.A0 (n_5866), .A1 (n_5864), .B0 (n_9931), .Y (n_9920));
AND2X1 g45909(.A (n_808), .B (n_528), .Y (n_12636));
NAND4X1 g45908(.A (n_4129), .B (n_4240), .C (n_1807), .D (n_1527), .Y(n_12635));
BUFX3 g40784(.A (n_937), .Y (n_4491));
NOR2X1 g40368(.A (n_2135), .B (n_2804), .Y (n_1937));
NOR2X1 g40369(.A (n_2006), .B (n_2684), .Y (n_1936));
NOR2X1 g40366(.A (n_2696), .B (n_2684), .Y (n_2650));
NOR2X1 g40367(.A (n_945), .B (n_2818), .Y (n_1938));
NOR2X1 g40364(.A (n_2470), .B (n_2712), .Y (n_1940));
NOR2X1 g40365(.A (n_867), .B (n_2831), .Y (n_1939));
NOR2X1 g40362(.A (n_2096), .B (n_2712), .Y (n_1941));
NOR2X1 g40363(.A (n_1016), .B (n_2712), .Y (n_2651));
AOI21X1 g40360(.A0 (oc5_cfg_1014), .A1 (in_slt_747), .B0(u14_u5_full_empty_r), .Y (n_554));
NOR2X1 g40361(.A (n_2749), .B (n_2716), .Y (n_2652));
NAND4X1 g37029(.A (n_2969), .B (n_3124), .C (n_1809), .D (n_1528), .Y(n_5818));
NAND4X1 g37028(.A (n_4131), .B (n_2281), .C (n_3188), .D (n_1545), .Y(n_6216));
AOI21X1 g38039(.A0 (u7_mem_b2_b_51 ), .A1 (n_4540), .B0 (n_1967), .Y(n_4516));
AOI21X1 g38038(.A0 (u3_mem_b2_b_36 ), .A1 (n_4519), .B0 (n_2032), .Y(n_4517));
AOI21X1 g38035(.A0 (u3_mem_b2_b_56 ), .A1 (n_4533), .B0 (n_2195), .Y(n_4521));
INVX1 g37022(.A (n_11855), .Y (n_5696));
NAND4X1 g37021(.A (n_4199), .B (n_3378), .C (n_2971), .D (n_1354), .Y(n_6202));
INVX1 g37020(.A (n_6202), .Y (n_5697));
INVX1 g37027(.A (n_6216), .Y (n_5692));
NAND4X1 g37026(.A (n_4190), .B (n_3171), .C (n_3848), .D (n_1529), .Y(n_5694));
INVX2 g37025(.A (n_5694), .Y (n_5693));
AOI21X1 g38032(.A0 (u6_mem_b2_b_47 ), .A1 (n_4544), .B0 (n_2319), .Y(n_4523));
NAND2X1 g36378(.A (n_6182), .B (n_2567), .Y (n_6292));
MX2X1 g38660(.A (u5_mem_b0_b_114 ), .B (wb_din_684), .S0 (n_3720), .Y(n_3714));
NAND2X1 g36370(.A (n_6216), .B (n_12634), .Y (n_6298));
NAND2X1 g36371(.A (n_6211), .B (n_12634), .Y (n_6297));
NAND2X1 g36372(.A (n_6233), .B (n_12634), .Y (n_6296));
NAND2X1 g36373(.A (n_6209), .B (n_12634), .Y (n_6295));
NAND2X1 g36376(.A (n_12514), .B (n_12634), .Y (n_6293));
NAND2X1 g36377(.A (n_5541), .B (n_12634), .Y (n_5914));
AOI22X1 g37769(.A0 (n_1756), .A1 (n_6368), .B0 (n_6515), .B1(n_1643), .Y (n_1666));
AND2X1 g30798(.A (n_9841), .B (n_11564), .Y (n_10394));
AOI21X1 g30799(.A0 (n_11948), .A1 (n_11949), .B0 (n_10945), .Y(n_10935));
AOI21X1 g30790(.A0 (n_12008), .A1 (n_12009), .B0 (n_10945), .Y(n_10947));
AOI21X1 g30791(.A0 (n_11988), .A1 (n_11989), .B0 (n_10945), .Y(n_10946));
AOI21X1 g30792(.A0 (n_12010), .A1 (n_12011), .B0 (n_10940), .Y(n_10944));
AOI21X1 g30793(.A0 (n_11674), .A1 (n_11675), .B0 (n_1473), .Y(n_10943));
AOI21X1 g30794(.A0 (n_11676), .A1 (n_11677), .B0 (n_1473), .Y(n_10942));
AOI21X1 g30795(.A0 (n_12000), .A1 (n_12001), .B0 (n_10940), .Y(n_10941));
AOI21X1 g30796(.A0 (n_11984), .A1 (n_11985), .B0 (n_1473), .Y(n_10939));
AOI21X1 g30797(.A0 (n_12018), .A1 (n_12019), .B0 (n_1473), .Y(n_10937));
NAND2X1 g38936(.A (u7_mem_b3_b_151 ), .B (n_1546), .Y (n_1522));
AOI22X1 g37689(.A0 (n_2558), .A1 (n_6390), .B0 (n_6660), .B1(n_2544), .Y (n_1695));
NAND2X1 g37688(.A (n_4136), .B (n_3036), .Y (n_5220));
NAND2X1 g37687(.A (n_4155), .B (n_2926), .Y (n_12851));
AOI21X1 g37685(.A0 (n_2558), .A1 (n_6375), .B0 (n_2257), .Y (n_3930));
NAND2X1 g37684(.A (n_4218), .B (n_2950), .Y (n_5222));
NAND2X1 g37683(.A (n_2607), .B (n_3401), .Y (n_4609));
AOI22X1 g37682(.A0 (n_6662), .A1 (n_2553), .B0 (n_6588), .B1(n_1316), .Y (n_2563));
NAND2X1 g37681(.A (n_2411), .B (n_3283), .Y (n_4610));
NAND2X1 g37680(.A (n_4112), .B (n_3490), .Y (n_12849));
INVX1 g41368(.A (n_1064), .Y (n_1851));
MX2X1 g31357(.A (u9_din_tmp_56), .B (in_slt_415), .S0 (n_9777), .Y(n_9780));
MX2X1 g31356(.A (u9_din_tmp_55), .B (in_slt_414), .S0 (n_9777), .Y(n_9782));
MX2X1 g31355(.A (u9_din_tmp_54), .B (in_slt_413), .S0 (n_9777), .Y(n_9784));
MX2X1 g31354(.A (u9_din_tmp_53), .B (in_slt_412), .S0 (n_9777), .Y(n_9785));
MX2X1 g31353(.A (u9_din_tmp_52), .B (in_slt_411), .S0 (n_9777), .Y(n_9786));
MX2X1 g31352(.A (u9_din_tmp_51), .B (in_slt_410), .S0 (n_9777), .Y(n_9788));
MX2X1 g31351(.A (u9_din_tmp1), .B (in_slt_400), .S0 (n_9777), .Y(n_9789));
MX2X1 g31350(.A (u10_din_tmp_46), .B (in_slt_427), .S0 (n_9860), .Y(n_9868));
MX2X1 g31359(.A (u9_din_tmp_43), .B (in_slt_402), .S0 (n_9777), .Y(n_9778));
MX2X1 g31358(.A (u9_din_tmp_42), .B (in_slt_401), .S0 (n_9777), .Y(n_9779));
NAND2X1 g31689(.A (n_288), .B (n_10391), .Y (n_10372));
NAND2X1 g31688(.A (n_129), .B (n_10391), .Y (n_10373));
NAND2X1 g31681(.A (n_1609), .B (n_10385), .Y (n_10382));
NAND2X1 g31680(.A (n_1614), .B (n_10391), .Y (n_10383));
NAND2X1 g31683(.A (n_1599), .B (n_10385), .Y (n_10379));
NAND2X1 g31682(.A (n_1604), .B (n_10376), .Y (n_10380));
NAND2X1 g31684(.A (n_1595), .B (n_10376), .Y (n_10378));
NAND2X1 g31687(.A (n_1580), .B (n_10385), .Y (n_10374));
NAND2X1 g31686(.A (n_1584), .B (n_10385), .Y (n_10375));
NAND2X1 g37979(.A (n_3213), .B (n_3524), .Y (n_5166));
NAND2X1 g37978(.A (n_2441), .B (n_2913), .Y (n_5167));
NAND2X1 g37971(.A (n_2410), .B (n_1915), .Y (n_4551));
NAND2X1 g34362(.A (u4_mem_b1_b_60 ), .B (n_7984), .Y (n_8041));
AOI22X1 g37973(.A0 (n_2502), .A1 (n_2500), .B0 (n_2499), .B1(n_1835), .Y (n_2501));
NAND2X1 g37972(.A (n_3158), .B (n_2974), .Y (n_5172));
NAND2X1 g37974(.A (n_2469), .B (n_3866), .Y (n_5171));
NAND2X1 g37977(.A (n_3411), .B (n_3082), .Y (n_5168));
NAND2X1 g37976(.A (n_3074), .B (n_3066), .Y (n_5169));
MX2X1 g36082(.A (n_6503), .B (n_6459), .S0 (n_6502), .Y (n_6504));
MX2X1 g36083(.A (n_5990), .B (n_5993), .S0 (n_6502), .Y (n_5991));
XOR2X1 g36080(.A (u26_ps_cnt_b3_b ), .B (n_1104), .Y (n_2630));
MX2X1 g36081(.A (n_6637), .B (n_6505), .S0 (n_6908), .Y (n_6506));
MX2X1 g36086(.A (n_6500), .B (n_6453), .S0 (n_6502), .Y (n_6501));
MX2X1 g36087(.A (n_6498), .B (n_6497), .S0 (n_6502), .Y (n_6499));
MX2X1 g36084(.A (n_5988), .B (n_5987), .S0 (n_6502), .Y (n_5989));
AND2X1 g33261(.A (n_5633), .B (u2_sync_resume), .Y (n_6067));
AOI21X1 g33260(.A0 (n_7458), .A1 (n_4730), .B0 (n_7353), .Y (n_8485));
NAND3X1 g33263(.A (n_862), .B (n_6838), .C (n_8101), .Y (n_8181));
NAND3X1 g33262(.A (n_8182), .B (u8_wp_b1_b ), .C (n_7976), .Y(n_8183));
NAND2X1 g41105(.A (oc3_cfg_995), .B (n_471), .Y (n_834));
AND2X1 g33264(.A (n_7521), .B (wb_din), .Y (n_7523));
NOR2X1 g41106(.A (wb_addr_i_b6_b), .B (n_593), .Y (n_594));
AOI22X1 g37880(.A0 (u11_din_tmp1), .A1 (n_4560), .B0 (n_4097), .B1(in_slt_442), .Y (n_3908));
INVX1 g45917(.A (n_12654), .Y (n_12656));
NOR2X1 g39979(.A (n_2218), .B (n_2767), .Y (n_2223));
NOR2X1 g39978(.A (n_2836), .B (n_2831), .Y (n_2840));
NAND2X1 g39973(.A (n_2325), .B (in_slt_452), .Y (n_1564));
NAND2X1 g39972(.A (n_11798), .B (u8_mem_b0_b_99 ), .Y (n_11449));
NAND2X1 g39971(.A (n_2491), .B (u7_mem_b0_b_115 ), .Y (n_1565));
NOR2X1 g39977(.A (n_945), .B (n_2732), .Y (n_2224));
NAND2X1 g38975(.A (u8_mem_b3_b_138 ), .B (n_2468), .Y (n_2386));
NOR2X1 g39975(.A (n_867), .B (n_2681), .Y (n_1838));
NAND2X1 g39974(.A (u8_mem_b1_b_87 ), .B (n_12291), .Y (n_2841));
NAND2X1 g45556(.A (n_12204), .B (u6_mem_b0_b_100 ), .Y (n_12164));
INVX2 g45915(.A (n_12659), .Y (n_12650));
NAND4X1 g45555(.A (n_12164), .B (n_12165), .C (n_12166), .D(n_12170), .Y (n_12171));
CLKBUFX3 g45550(.A (n_12503), .Y (n_12161));
AOI22X1 g37885(.A0 (u10_din_tmp_56), .A1 (n_3339), .B0 (n_3911), .B1(in_slt_435), .Y (n_3904));
NAND2X1 g34831(.A (u8_mem_b1_b_81 ), .B (n_7976), .Y (n_7603));
NAND2X1 g34830(.A (u8_mem_b1_b_80 ), .B (n_7976), .Y (n_7604));
NAND2X1 g34833(.A (u8_mem_b1_b_84 ), .B (n_7976), .Y (n_7601));
NAND2X1 g34832(.A (u8_mem_b1_b_83 ), .B (n_7976), .Y (n_7602));
NAND2X1 g34835(.A (u8_mem_b1_b_85 ), .B (n_7976), .Y (n_7599));
NAND2X1 g34834(.A (u3_mem_b1_b ), .B (n_8141), .Y (n_7600));
NAND2X1 g34837(.A (u3_mem_b1_b_69 ), .B (n_8101), .Y (n_7597));
NAND2X1 g34836(.A (u8_mem_b1_b_86 ), .B (n_7976), .Y (n_7598));
NAND2X1 g34838(.A (u8_mem_b1_b_87 ), .B (n_7976), .Y (n_7596));
AOI21X1 g38314(.A0 (u5_mem_b2_b_29 ), .A1 (n_4370), .B0 (n_2114), .Y(n_4368));
XOR2X1 g35496(.A (n_5620), .B (n_4092), .Y (n_5621));
AOI22X1 g37884(.A0 (u11_din_tmp_52), .A1 (n_4560), .B0 (n_4097), .B1(in_slt_453), .Y (n_3905));
NOR2X1 g35300(.A (n_1301), .B (n_12335), .Y (n_7542));
OR2X1 g35301(.A (n_5831), .B (n_11827), .Y (n_8669));
INVX1 g35302(.A (n_8667), .Y (n_9478));
INVX1 g35303(.A (n_7541), .Y (n_8667));
NOR2X1 g35304(.A (n_1372), .B (n_12335), .Y (n_7541));
OR2X1 g35305(.A (n_2485), .B (n_11827), .Y (n_8666));
INVX1 g35306(.A (n_8665), .Y (n_9477));
INVX1 g35307(.A (n_7539), .Y (n_8665));
OR2X1 g35309(.A (n_5827), .B (n_11827), .Y (n_8664));
NAND2X1 g39355(.A (u8_mem_b2_b_29 ), .B (n_3334), .Y (n_11741));
NAND2X1 g39354(.A (u5_mem_b2_b_39 ), .B (n_12823), .Y (n_12033));
NAND2X1 g39353(.A (n_3259), .B (u5_mem_b0_b_101 ), .Y (n_3251));
NAND2X1 g39352(.A (n_3252), .B (u7_mem_b0_b_120 ), .Y (n_3253));
NAND2X1 g39351(.A (n_3259), .B (u5_mem_b0_b_99 ), .Y (n_3254));
NAND2X1 g39350(.A (u5_mem_b2_b_51 ), .B (n_12823), .Y (n_2320));
NAND4X1 g36969(.A (n_11713), .B (n_11714), .C (n_2482), .D (n_1869),.Y (n_5835));
INVX1 g36968(.A (n_5835), .Y (n_5555));
NAND4X1 g36965(.A (n_11751), .B (n_11752), .C (n_2229), .D (n_2431),.Y (n_5844));
INVX1 g36964(.A (n_5844), .Y (n_5556));
NAND4X1 g36967(.A (n_11670), .B (n_11671), .C (n_1786), .D (n_4250),.Y (n_6805));
INVX1 g36966(.A (n_6805), .Y (n_6077));
NAND2X1 g36961(.A (n_1586), .B (n_1583), .Y (n_4008));
NAND2X1 g36960(.A (n_1588), .B (n_1587), .Y (n_4009));
NAND2X1 g36963(.A (n_1579), .B (n_1578), .Y (n_4006));
AOI21X1 g38334(.A0 (u5_mem_b2_b_36 ), .A1 (n_4370), .B0 (n_2476), .Y(n_4352));
AOI22X1 g37886(.A0 (u11_din_tmp_53), .A1 (n_4560), .B0 (n_4097), .B1(in_slt_454), .Y (n_3903));
INVX4 g45911(.A (n_12636), .Y (n_12640));
AOI21X1 g38335(.A0 (u6_mem_b1_b_80 ), .A1 (n_5019), .B0 (n_2660), .Y(n_5003));
NAND2X1 g31(.A (n_12355), .B (n_12358), .Y (n_12359));
AOI21X1 g30(.A0 (u4_mem_b0_b_105 ), .A1 (n_12840), .B0 (n_11842), .Y(n_11843));
NAND2X2 g33(.A (n_761), .B (n_445), .Y (n_11844));
NAND2X1 g32(.A (n_12746), .B (n_12357), .Y (n_12358));
INVX4 g35(.A (n_11851), .Y (n_11852));
AND2X1 g34(.A (n_12087), .B (u4_mem_b2_b_43 ), .Y (n_11842));
AND2X1 g37(.A (n_283), .B (oc1_cfg_975), .Y (n_12357));
INVX2 g36(.A (n_12333), .Y (n_11851));
NAND2X1 g39(.A (n_12261), .B (u4_mem_b1_b_72 ), .Y (n_12740));
OAI21X1 g38(.A0 (n_5687), .A1 (n_7088), .B0 (n_6146), .Y (n_12125));
INVX4 g40462(.A (wb_din_664), .Y (n_2794));
INVX2 g40469(.A (wb_din_679), .Y (n_2818));
NAND2X1 g34309(.A (u3_mem_b3_b_143 ), .B (n_8101), .Y (n_8087));
NAND2X1 g34308(.A (u3_mem_b3_b_142 ), .B (n_8101), .Y (n_8088));
OAI21X1 g33467(.A0 (n_4512), .A1 (n_8440), .B0 (n_8107), .Y (n_8392));
NAND2X1 g34306(.A (n_6706), .B (n_7475), .Y (n_8245));
OAI21X1 g33465(.A0 (n_4324), .A1 (n_8911), .B0 (n_8110), .Y (n_8395));
OAI21X1 g33464(.A0 (n_4293), .A1 (n_8856), .B0 (n_8112), .Y (n_8396));
OAI21X1 g33463(.A0 (n_4394), .A1 (n_8097), .B0 (n_8113), .Y (n_8397));
OAI21X1 g33462(.A0 (n_4480), .A1 (n_8097), .B0 (n_8114), .Y (n_8398));
NAND2X1 g34301(.A (u3_mem_b3_b_137 ), .B (n_8097), .Y (n_8094));
OAI21X1 g33460(.A0 (n_4518), .A1 (n_8097), .B0 (n_8116), .Y (n_8400));
AOI21X1 g38484(.A0 (u7_mem_b1_b_84 ), .A1 (n_5069), .B0 (n_2840), .Y(n_4896));
AOI21X1 g38485(.A0 (u7_mem_b1_b_86 ), .A1 (n_5069), .B0 (n_2656), .Y(n_4895));
AOI21X1 g38486(.A0 (u7_mem_b1_b_88 ), .A1 (n_5069), .B0 (n_2715), .Y(n_4894));
AOI21X1 g38487(.A0 (u7_mem_b1_b_89 ), .A1 (n_5069), .B0 (n_2647), .Y(n_4893));
AOI21X1 g38480(.A0 (u7_mem_b1_b_76 ), .A1 (n_5118), .B0 (n_2706), .Y(n_4900));
AOI21X1 g38481(.A0 (u7_mem_b1_b_80 ), .A1 (n_5069), .B0 (n_2730), .Y(n_4899));
AOI21X1 g38482(.A0 (u7_mem_b3_b_145 ), .A1 (n_5145), .B0 (n_3103), .Y(n_4898));
AOI21X1 g38483(.A0 (u7_mem_b1_b_82 ), .A1 (n_5069), .B0 (n_2649), .Y(n_4897));
AOI21X1 g38488(.A0 (u7_mem_b1_b_62 ), .A1 (n_5118), .B0 (n_2805), .Y(n_4892));
AOI21X1 g38489(.A0 (u7_mem_b1_b_66 ), .A1 (n_5069), .B0 (n_2714), .Y(n_4891));
INVX1 g40879(.A (n_1430), .Y (n_2751));
NAND2X1 g39321(.A (u3_mem_b2_b_33 ), .B (n_12619), .Y (n_11738));
AOI21X1 g38260(.A0 (u6_mem_b3_b_141 ), .A1 (n_5059), .B0 (n_3177), .Y(n_5051));
AOI21X1 g38261(.A0 (u6_mem_b3_b_122 ), .A1 (n_5100), .B0 (n_3164), .Y(n_5050));
AOI21X1 g38262(.A0 (u5_mem_b1_b ), .A1 (n_5048), .B0 (n_2802), .Y(n_5049));
AOI21X1 g38263(.A0 (u5_mem_b1_b_69 ), .A1 (n_5048), .B0 (n_2760), .Y(n_5047));
AOI21X1 g38264(.A0 (u5_mem_b1_b_70 ), .A1 (n_5048), .B0 (n_2717), .Y(n_5046));
AOI21X1 g38265(.A0 (u3_mem_b3_b_141 ), .A1 (n_5133), .B0 (n_3428), .Y(n_5045));
AOI21X1 g38266(.A0 (u6_mem_b3_b_139 ), .A1 (n_5059), .B0 (n_3344), .Y(n_5044));
AOI21X1 g38267(.A0 (u8_mem_b1_b_77 ), .A1 (n_4387), .B0 (n_2051), .Y(n_4383));
AOI21X1 g38268(.A0 (u5_mem_b1_b_72 ), .A1 (n_5048), .B0 (n_2725), .Y(n_5043));
AOI21X1 g38269(.A0 (u5_mem_b1_b_73 ), .A1 (n_5048), .B0 (n_2785), .Y(n_5042));
AOI22X1 g37767(.A0 (n_2558), .A1 (n_6386), .B0 (n_6610), .B1(n_2534), .Y (n_2535));
AOI22X1 g37760(.A0 (n_42), .A1 (n_2553), .B0 (n_5510), .B1 (n_1316),.Y (n_2537));
AOI22X1 g37761(.A0 (n_1756), .A1 (n_6377), .B0 (n_6522), .B1(n_1643), .Y (n_1672));
AOI22X1 g37762(.A0 (n_6526), .A1 (n_2530), .B0 (n_6652), .B1(n_2534), .Y (n_2536));
AOI21X1 g37763(.A0 (n_6554), .A1 (n_1831), .B0 (n_1215), .Y (n_1671));
NAND2X1 g39326(.A (u5_mem_b1_b_87 ), .B (n_3209), .Y (n_3274));
OAI21X1 g33078(.A0 (n_7209), .A1 (n_7056), .B0 (n_10481), .Y(n_11735));
OAI21X1 g33079(.A0 (n_7117), .A1 (n_6978), .B0 (n_10483), .Y(n_11629));
OAI21X1 g33074(.A0 (n_7118), .A1 (n_6979), .B0 (n_10483), .Y(n_11623));
OAI21X1 g33075(.A0 (n_7211), .A1 (n_7059), .B0 (n_12689), .Y(n_11731));
OAI21X1 g33076(.A0 (n_7210), .A1 (n_7058), .B0 (n_12689), .Y(n_11733));
OAI21X1 g33077(.A0 (n_7124), .A1 (n_7057), .B0 (n_10483), .Y(n_11625));
OAI21X1 g33070(.A0 (n_7215), .A1 (n_7062), .B0 (n_10481), .Y(n_12062));
OAI21X1 g33071(.A0 (n_7119), .A1 (n_6982), .B0 (n_10483), .Y(n_11627));
OAI21X1 g33072(.A0 (n_7244), .A1 (n_11901), .B0 (n_10481), .Y(n_11994));
OAI21X1 g33073(.A0 (n_7213), .A1 (n_7060), .B0 (n_10483), .Y(n_11621));
NOR2X1 g37508(.A (n_4751), .B (n_6594), .Y (n_3956));
NAND2X1 g39420(.A (u4_mem_b1_b_60 ), .B (n_12272), .Y (n_4195));
NAND2X1 g39423(.A (n_4560), .B (in_slt_458), .Y (n_5296));
NAND2X1 g39327(.A (u8_mem_b1_b_61 ), .B (n_12291), .Y (n_12843));
AND2X1 g30911(.A (n_9960), .B (n_11600), .Y (n_10778));
NAND2X1 g39425(.A (u5_mem_b1_b_64 ), .B (n_3257), .Y (n_12809));
MX2X1 g38689(.A (u6_mem_b0_b_92 ), .B (wb_din_662), .S0 (n_3632), .Y(n_3668));
NAND2X1 g39424(.A (u8_mem_b1_b_79 ), .B (n_12291), .Y (n_3191));
NOR2X1 g39427(.A (u11_mem_b2_b_98 ), .B (n_1214), .Y (n_1005));
NAND2X1 g39426(.A (n_2344), .B (in_slt_423), .Y (n_2305));
OAI21X1 g33816(.A0 (n_5128), .A1 (n_9055), .B0 (n_7710), .Y (n_9052));
NAND2X1 g34265(.A (u3_mem_b2_b_41 ), .B (n_8101), .Y (n_8136));
OAI21X1 g33546(.A0 (n_4433), .A1 (n_8333), .B0 (n_8011), .Y (n_8294));
NOR2X1 g40194(.A (n_2720), .B (n_933), .Y (n_2051));
NOR2X1 g40197(.A (n_2477), .B (n_2702), .Y (n_2048));
NAND2X1 g34267(.A (u8_mem_b3_b_126 ), .B (n_7976), .Y (n_8133));
NOR2X1 g40191(.A (n_1082), .B (n_2735), .Y (n_2726));
NOR2X1 g40190(.A (n_2154), .B (n_2818), .Y (n_2319));
NOR2X1 g40193(.A (n_1082), .B (n_2681), .Y (n_2725));
NAND2X1 g40192(.A (n_5118), .B (n_4540), .Y (n_2052));
OAI21X1 g33540(.A0 (n_4441), .A1 (n_9349), .B0 (n_8017), .Y (n_8301));
NOR2X1 g40199(.A (n_2721), .B (n_2720), .Y (n_2722));
NOR2X1 g40198(.A (n_2470), .B (n_2744), .Y (n_2047));
OAI21X1 g33813(.A0 (n_5110), .A1 (n_9034), .B0 (n_7715), .Y (n_9058));
NAND2X1 g34611(.A (u6_mem_b1_b_79 ), .B (n_7758), .Y (n_7815));
OAI21X1 g33542(.A0 (n_4310), .A1 (n_8318), .B0 (n_8015), .Y (n_8298));
NAND2X1 g34610(.A (u6_mem_b1_b_60 ), .B (n_7758), .Y (n_7817));
OAI21X1 g33543(.A0 (n_4438), .A1 (n_9349), .B0 (n_8014), .Y (n_8297));
NAND2X1 g34613(.A (u6_mem_b1_b_81 ), .B (n_7758), .Y (n_7812));
NAND2X1 g34612(.A (u6_mem_b1_b_80 ), .B (n_7758), .Y (n_7813));
NAND2X1 g36419(.A (n_6260), .B (n_6259), .Y (n_6261));
MX2X1 g36149(.A (n_6845), .B (n_6906), .S0 (n_6856), .Y (n_6846));
MX2X1 g36148(.A (n_6394), .B (n_6560), .S0 (n_6856), .Y (n_6395));
MX2X1 g36147(.A (n_6847), .B (n_6927), .S0 (n_6856), .Y (n_6848));
NAND2X1 g34615(.A (u6_mem_b1_b_83 ), .B (n_7758), .Y (n_7810));
MX2X1 g36145(.A (n_6852), .B (n_6913), .S0 (n_6856), .Y (n_6853));
MX2X1 g36144(.A (n_6854), .B (n_6896), .S0 (n_6856), .Y (n_6855));
MX2X1 g36142(.A (n_6859), .B (n_6916), .S0 (n_6856), .Y (n_6860));
MX2X1 g36141(.A (n_6862), .B (n_6920), .S0 (n_6856), .Y (n_6863));
NAND2X1 g34614(.A (u6_mem_b1_b_82 ), .B (n_7758), .Y (n_7811));
INVX1 g42739(.A (n_458), .Y (n_991));
MX2X1 g36132(.A (n_5966), .B (n_6003), .S0 (n_6475), .Y (n_5967));
NAND2X1 g34617(.A (u6_mem_b1_b_85 ), .B (n_7758), .Y (n_7808));
OAI21X1 g33548(.A0 (n_4431), .A1 (n_8333), .B0 (n_8009), .Y (n_8291));
INVX1 g42731(.A (n_1473), .Y (n_2343));
NAND2X1 g34616(.A (u6_mem_b1_b_84 ), .B (n_7758), .Y (n_7809));
INVX2 g42737(.A (n_991), .Y (n_1473));
INVX1 g42735(.A (n_991), .Y (n_10945));
OAI21X1 g33549(.A0 (n_4430), .A1 (n_9333), .B0 (n_8008), .Y (n_8290));
NAND2X1 g34619(.A (u6_mem_b1_b_87 ), .B (n_7758), .Y (n_7806));
INVX1 g40998(.A (n_1416), .Y (n_2780));
NOR2X1 g37505(.A (n_4761), .B (n_6594), .Y (n_3958));
NAND2X1 g40994(.A (n_434), .B (n_4690), .Y (n_1156));
BUFX3 g40997(.A (n_1016), .Y (n_5148));
BUFX3 g40996(.A (n_1016), .Y (n_5157));
INVX4 g40992(.A (n_1156), .Y (n_2344));
NOR2X1 g35829(.A (n_5248), .B (n_5225), .Y (n_5226));
NOR2X1 g35828(.A (n_5248), .B (wb_addr_i_b6_b), .Y (n_6045));
INVX8 g41648(.A (n_1111), .Y (n_2468));
NOR2X1 g35821(.A (n_513), .B (n_6752), .Y (n_6755));
NOR2X1 g35820(.A (n_609), .B (n_6752), .Y (n_6754));
NOR2X1 g35823(.A (n_617), .B (n_6752), .Y (n_6759));
NOR2X1 g35822(.A (n_750), .B (n_6752), .Y (n_6758));
NOR2X1 g35825(.A (n_541), .B (n_5440), .Y (n_6062));
NOR2X1 g35824(.A (n_733), .B (n_6752), .Y (n_6671));
NOR2X1 g35827(.A (n_666), .B (n_6752), .Y (n_6064));
NOR2X1 g35826(.A (n_550), .B (n_5440), .Y (n_6063));
INVX1 g42597(.A (u10_mem_b3_b_57 ), .Y (n_6007));
INVX1 g42595(.A (u10_mem_b0_b_166 ), .Y (n_5955));
INVX1 g42594(.A (u10_mem_b3_b_72 ), .Y (n_6013));
INVX1 g42591(.A (u11_mem_b2_b_114 ), .Y (n_236));
INVX1 g42590(.A (u11_mem_b1_b_138 ), .Y (n_1633));
AOI21X1 g38034(.A0 (u5_mem_b1_b_67 ), .A1 (n_5048), .B0 (n_2774), .Y(n_5141));
INVX1 g42599(.A (n_763), .Y (n_814));
MX2X1 g36130(.A (n_6408), .B (n_6566), .S0 (n_6475), .Y (n_6409));
AOI22X1 g37660(.A0 (in_slt_412), .A1 (n_1406), .B0 (in_slt_414), .B1(n_4624), .Y (n_4626));
NAND2X1 g38933(.A (u7_mem_b3_b_135 ), .B (n_1538), .Y (n_1524));
INVX2 g40700(.A (n_1434), .Y (n_3441));
CLKBUFX1 g40821(.A (n_806), .Y (n_6995));
INVX1 g40702(.A (n_1178), .Y (n_1434));
INVX1 g40820(.A (n_6995), .Y (n_1229));
INVX1 g40704(.A (n_2366), .Y (n_1549));
NAND2X1 g39004(.A (u3_mem_b1_b_84 ), .B (n_3316), .Y (n_3521));
INVX1 g40822(.A (n_806), .Y (n_5881));
AOI21X1 g30817(.A0 (n_9925), .A1 (n_9806), .B0 (n_10916), .Y(n_10917));
AOI21X1 g30816(.A0 (n_9926), .A1 (n_9807), .B0 (n_2485), .Y(n_10919));
AOI21X1 g30815(.A0 (n_9927), .A1 (n_9808), .B0 (n_2485), .Y(n_10920));
AOI21X1 g30814(.A0 (n_9928), .A1 (n_9810), .B0 (n_10921), .Y(n_10922));
AOI21X1 g30813(.A0 (n_9929), .A1 (n_9811), .B0 (n_10916), .Y(n_10923));
AOI21X1 g30812(.A0 (n_9930), .A1 (n_9812), .B0 (n_10921), .Y(n_10924));
AOI21X1 g30811(.A0 (n_9932), .A1 (n_9813), .B0 (n_2485), .Y(n_10926));
AOI21X1 g30810(.A0 (n_9933), .A1 (n_9815), .B0 (n_2485), .Y(n_10927));
NOR2X1 g39508(.A (n_3117), .B (n_2735), .Y (n_3133));
NOR2X1 g39509(.A (n_3117), .B (n_2818), .Y (n_3132));
AOI22X1 g37662(.A0 (in_slt_415), .A1 (n_4623), .B0 (in_slt_403), .B1(n_2368), .Y (n_5733));
MX2X1 g31306(.A (n_5653), .B (n_1620), .S0 (n_9721), .Y (n_10441));
AOI21X1 g30819(.A0 (n_9922), .A1 (n_9804), .B0 (n_10921), .Y(n_10914));
AOI21X1 g30818(.A0 (n_12835), .A1 (n_12836), .B0 (n_2485), .Y(n_10915));
MX2X1 g34152(.A (u8_mem_b0_b_119 ), .B (n_3587), .S0 (n_7490), .Y(n_9376));
MX2X1 g34153(.A (u8_mem_b0_b_92 ), .B (n_3746), .S0 (n_7490), .Y(n_8693));
MX2X1 g34150(.A (u3_mem_b0_b_115 ), .B (n_3588), .S0 (n_8700), .Y(n_8694));
MX2X1 g31307(.A (n_5665), .B (n_1246), .S0 (n_10315), .Y (n_10130));
MX2X1 g34156(.A (u8_mem_b0_b_121 ), .B (n_3822), .S0 (n_7490), .Y(n_8692));
MX2X1 g34157(.A (u8_mem_b0_b_93 ), .B (n_3832), .S0 (n_7490), .Y(n_8691));
MX2X1 g34154(.A (u8_mem_b0_b_120 ), .B (n_3748), .S0 (n_7490), .Y(n_9375));
MX2X1 g34155(.A (u3_mem_b0_b_117 ), .B (n_3585), .S0 (n_8700), .Y(n_9373));
NAND2X1 g31652(.A (n_1732), .B (n_10045), .Y (n_9995));
MX2X1 g34158(.A (u8_mem_b0_b_94 ), .B (n_3837), .S0 (n_7490), .Y(n_9371));
MX2X1 g34159(.A (u8_mem_b0_b_95 ), .B (n_3583), .S0 (n_7490), .Y(n_9370));
MX2X1 g31301(.A (n_6389), .B (n_6388), .S0 (n_9818), .Y (n_10812));
AOI21X1 g38030(.A0 (u3_mem_b2_b_50 ), .A1 (n_4533), .B0 (n_2147), .Y(n_4524));
MX2X1 g31302(.A (n_5950), .B (n_5949), .S0 (n_10450), .Y (n_10446));
AOI22X1 g37665(.A0 (n_2502), .A1 (n_1704), .B0 (n_1703), .B1(n_1859), .Y (n_1705));
MX2X1 g31303(.A (n_5657), .B (n_1634), .S0 (n_10513), .Y (n_10445));
NAND2X1 g39002(.A (u7_mem_b1_b_79 ), .B (n_3522), .Y (n_3523));
NAND2X1 g39123(.A (u9_din_tmp_49), .B (n_2368), .Y (n_1925));
AOI22X1 g37664(.A0 (n_2558), .A1 (n_1251), .B0 (n_5506), .B1(n_1316), .Y (n_1252));
OR2X1 g41618(.A (n_469), .B (n_12584), .Y (n_977));
OAI21X1 g33898(.A0 (n_4957), .A1 (n_8948), .B0 (n_7625), .Y (n_8950));
OAI21X1 g33899(.A0 (n_4931), .A1 (n_8948), .B0 (n_7624), .Y (n_8949));
OAI21X1 g33896(.A0 (n_4912), .A1 (n_8951), .B0 (n_7627), .Y (n_8953));
OAI21X1 g33897(.A0 (n_4878), .A1 (n_8951), .B0 (n_7626), .Y (n_8952));
OAI21X1 g33894(.A0 (n_4909), .A1 (n_8961), .B0 (n_7630), .Y (n_8955));
OAI21X1 g33895(.A0 (n_4879), .A1 (n_8961), .B0 (n_7628), .Y (n_8954));
OAI21X1 g33892(.A0 (n_4876), .A1 (n_8958), .B0 (n_7632), .Y (n_8957));
OAI21X1 g33893(.A0 (n_4880), .A1 (n_8958), .B0 (n_7631), .Y (n_8956));
OAI21X1 g33890(.A0 (n_4862), .A1 (n_8958), .B0 (n_7634), .Y (n_8960));
OAI21X1 g33891(.A0 (n_4959), .A1 (n_8958), .B0 (n_7633), .Y (n_8959));
AOI22X1 g37667(.A0 (in_slt_399), .A1 (n_4623), .B0 (u9_din_tmp_44),.B1 (n_4616), .Y (n_4618));
MX2X1 g38729(.A (u7_mem_b0_b_92 ), .B (wb_din_662), .S0 (n_3622), .Y(n_3612));
NOR2X1 g39000(.A (n_3486), .B (n_2744), .Y (n_3525));
AOI21X1 g38098(.A0 (u3_mem_b2_b_59 ), .A1 (n_4533), .B0 (n_2108), .Y(n_4480));
NOR2X1 g39125(.A (n_2790), .B (n_1488), .Y (n_1496));
AOI21X1 g38097(.A0 (u7_mem_b2_b_52 ), .A1 (n_4540), .B0 (n_2104), .Y(n_4481));
AOI21X1 g38096(.A0 (u3_mem_b3_b_145 ), .A1 (n_5138), .B0 (n_2947), .Y(n_5120));
NOR2X1 g37511(.A (n_5339), .B (n_6594), .Y (n_4655));
NOR2X1 g37510(.A (n_5330), .B (n_6594), .Y (n_4656));
NAND2X1 g39507(.A (n_12389), .B (u4_mem_b0_b_115 ), .Y (n_3134));
MX2X1 g38721(.A (u6_mem_b0_b_118 ), .B (wb_din_688), .S0 (n_3632), .Y(n_3621));
INVX1 g37040(.A (n_6207), .Y (n_5688));
NOR2X1 g37515(.A (n_5315), .B (n_6649), .Y (n_4654));
AOI21X1 g38090(.A0 (u3_mem_b2_b_45 ), .A1 (n_4533), .B0 (n_2072), .Y(n_4484));
NOR2X1 g40205(.A (n_2780), .B (n_2801), .Y (n_3412));
NOR2X1 g40204(.A (n_2043), .B (n_2801), .Y (n_2044));
NOR2X1 g40207(.A (n_2041), .B (n_2735), .Y (n_2042));
NOR2X1 g40206(.A (n_2748), .B (n_2067), .Y (n_2351));
NOR2X1 g40201(.A (n_1016), .B (n_2794), .Y (n_2718));
NOR2X1 g40200(.A (n_2759), .B (n_2748), .Y (n_2719));
NOR2X1 g40203(.A (n_2712), .B (n_2045), .Y (n_2046));
NOR2X1 g40202(.A (n_2784), .B (n_2716), .Y (n_2717));
NAND2X1 g39127(.A (in_slt_400), .B (n_2368), .Y (n_2354));
AOI21X1 g40208(.A0 (oc4_cfg_1004), .A1 (in_slt_748), .B0(u14_u4_full_empty_r), .Y (n_539));
NAND2X1 g39582(.A (u6_mem_b1_b_71 ), .B (n_12169), .Y (n_4164));
INVX1 g43058(.A (u10_mem_b0_b_167 ), .Y (n_314));
AND2X1 g45927(.A (n_925), .B (oc0_cfg_965), .Y (n_12664));
NAND2X1 g45926(.A (n_12664), .B (n_12755), .Y (n_12666));
AOI22X1 g37742(.A0 (n_2558), .A1 (n_1240), .B0 (n_5357), .B1(n_1316), .Y (n_1241));
AOI21X1 g45924(.A0 (n_6289), .A1 (n_5762), .B0 (n_7214), .Y(n_12663));
OAI21X1 g45923(.A0 (n_12663), .A1 (n_12668), .B0 (n_10481), .Y(n_12672));
INVX2 g45922(.A (n_12509), .Y (n_12662));
INVX2 g45921(.A (n_12662), .Y (n_12659));
AOI21X1 g38017(.A0 (u3_mem_b2_b_40 ), .A1 (n_4533), .B0 (n_2127), .Y(n_4532));
AOI21X1 g38015(.A0 (u6_mem_b2_b_50 ), .A1 (n_4544), .B0 (n_2186), .Y(n_4535));
AOI21X1 g38014(.A0 (u8_mem_b3_b_149 ), .A1 (n_3879), .B0 (n_1283), .Y(n_3887));
AOI21X1 g38013(.A0 (u7_mem_b2_b_57 ), .A1 (n_4540), .B0 (n_2217), .Y(n_4536));
AOI21X1 g38012(.A0 (u3_mem_b2_b ), .A1 (n_4533), .B0 (n_2105), .Y(n_4537));
AOI21X1 g38011(.A0 (u3_mem_b1_b_68 ), .A1 (n_5148), .B0 (n_2678), .Y(n_5147));
AOI21X1 g38010(.A0 (u7_mem_b2_b_30 ), .A1 (n_4540), .B0 (n_2203), .Y(n_4538));
NOR2X1 g40340(.A (n_2144), .B (n_3008), .Y (n_1953));
NOR2X1 g40341(.A (n_2189), .B (n_2681), .Y (n_1952));
NOR2X1 g40342(.A (n_867), .B (n_2767), .Y (n_1951));
NOR2X1 g40343(.A (n_2085), .B (n_2794), .Y (n_1950));
NOR2X1 g40344(.A (n_2749), .B (n_2686), .Y (n_2659));
NOR2X1 g40345(.A (n_867), .B (n_2763), .Y (n_1949));
AOI21X1 g38019(.A0 (u8_mem_b2_b_37 ), .A1 (n_4499), .B0 (n_2196), .Y(n_4530));
AOI21X1 g38018(.A0 (u6_mem_b2_b_49 ), .A1 (n_4544), .B0 (n_1800), .Y(n_4531));
NAND2X1 g37743(.A (n_1328), .B (n_4171), .Y (n_5214));
INVX1 g43053(.A (u9_mem_b2_b_110 ), .Y (n_1561));
NAND2X1 g39580(.A (u8_mem_b2_b_57 ), .B (n_3441), .Y (n_3084));
NAND2X1 g37740(.A (n_3069), .B (n_3846), .Y (n_4598));
AOI21X1 g38095(.A0 (u8_mem_b2_b_58 ), .A1 (n_4491), .B0 (n_2159), .Y(n_4482));
AOI22X1 g37741(.A0 (n_2502), .A1 (n_6852), .B0 (n_6945), .B1(n_1859), .Y (n_1674));
AOI21X1 g38094(.A0 (u8_mem_b2_b_59 ), .A1 (n_4499), .B0 (n_1982), .Y(n_4483));
INVX1 g42769(.A (u11_mem_b2_b_108 ), .Y (n_1627));
NAND2X1 g39587(.A (u6_mem_b2_b_53 ), .B (n_3423), .Y (n_3080));
INVX4 g41347(.A (n_1134), .Y (n_5371));
XOR2X1 g38093(.A (u11_rp_b2_b ), .B (n_736), .Y (n_1080));
OAI21X1 g33799(.A0 (n_5058), .A1 (n_9077), .B0 (n_7728), .Y (n_9073));
OAI21X1 g33798(.A0 (n_4914), .A1 (n_9077), .B0 (n_7729), .Y (n_9074));
OR2X1 g36310(.A (n_2621), .B (n_3942), .Y (n_2622));
NAND2X1 g36311(.A (n_6161), .B (n_6316), .Y (n_6325));
NAND2X1 g36316(.A (n_12354), .B (n_6824), .Y (n_6833));
NAND2X1 g36314(.A (n_6244), .B (n_2567), .Y (n_6324));
NAND2X1 g36315(.A (n_6777), .B (n_6824), .Y (n_6834));
OAI21X1 g33791(.A0 (n_5062), .A1 (n_9105), .B0 (n_7736), .Y (n_9083));
OAI21X1 g33790(.A0 (n_4919), .A1 (n_9105), .B0 (n_7737), .Y (n_9084));
OAI21X1 g33793(.A0 (n_5109), .A1 (n_9080), .B0 (n_7734), .Y (n_9081));
OAI21X1 g33794(.A0 (n_4917), .A1 (n_9077), .B0 (n_7733), .Y (n_9079));
OAI21X1 g33797(.A0 (n_4915), .A1 (n_9080), .B0 (n_7730), .Y (n_9075));
OAI21X1 g33796(.A0 (n_4916), .A1 (n_9080), .B0 (n_7731), .Y (n_9076));
MX2X1 g31331(.A (n_5469), .B (n_1238), .S0 (n_9724), .Y (n_10418));
MX2X1 g31330(.A (n_6350), .B (n_6349), .S0 (n_10537), .Y (n_10420));
MX2X1 g31333(.A (n_6345), .B (n_6344), .S0 (n_10537), .Y (n_10416));
MX2X1 g31335(.A (n_5948), .B (n_5947), .S0 (n_10537), .Y (n_10413));
MX2X1 g31334(.A (n_5639), .B (n_2539), .S0 (n_10565), .Y (n_10415));
MX2X1 g31337(.A (n_5643), .B (n_1251), .S0 (n_10315), .Y (n_10127));
MX2X1 g31336(.A (n_6343), .B (n_6342), .S0 (n_10565), .Y (n_10412));
MX2X1 g31339(.A (n_6340), .B (n_6339), .S0 (n_10315), .Y (n_10124));
MX2X1 g31338(.A (n_5641), .B (n_1864), .S0 (n_10315), .Y (n_10126));
INVX2 g40838(.A (n_867), .Y (n_1167));
INVX1 g40839(.A (n_1167), .Y (n_2171));
OAI21X1 g37405(.A0 (u10_mem_b0_b_175 ), .A1 (n_6341), .B0 (n_4641), .Y(n_5471));
OAI21X1 g37404(.A0 (u10_mem_b0_b_174 ), .A1 (n_5645), .B0 (n_5230), .Y(n_5646));
OAI21X1 g37407(.A0 (u10_mem_b0_b_177 ), .A1 (n_6341), .B0 (n_4653), .Y(n_5469));
OAI21X1 g37406(.A0 (u10_mem_b0_b_176 ), .A1 (n_6341), .B0 (n_4648), .Y(n_5470));
OAI21X1 g37401(.A0 (u10_mem_b0_b_172 ), .A1 (n_6341), .B0 (n_5232), .Y(n_5649));
OAI21X1 g37400(.A0 (u11_mem_b0_b_175 ), .A1 (n_6359), .B0 (n_5237), .Y(n_5650));
OAI21X1 g37403(.A0 (u10_mem_b0_b_173 ), .A1 (n_5645), .B0 (n_5231), .Y(n_5647));
OAI21X1 g37402(.A0 (u11_mem_b0_b_179 ), .A1 (n_6359), .B0 (n_5243), .Y(n_5648));
NAND2X1 g37959(.A (n_2456), .B (n_2896), .Y (n_5181));
NAND2X1 g37958(.A (n_3862), .B (n_3136), .Y (n_5182));
OAI21X1 g37408(.A0 (u11_mem_b0_b_177 ), .A1 (n_6359), .B0 (n_5234), .Y(n_5644));
XOR2X1 g38091(.A (u9_wp_b3_b ), .B (n_1063), .Y (n_3875));
INVX1 g33249(.A (u15_crac_we_r), .Y (n_8486));
NAND2X1 g37745(.A (n_2401), .B (n_2317), .Y (n_3915));
AOI21X1 g38355(.A0 (u5_mem_b3_b_145 ), .A1 (n_4996), .B0 (n_3128), .Y(n_4982));
NAND2X1 g36392(.A (n_5807), .B (n_2567), .Y (n_5908));
NAND2X1 g34305(.A (u3_mem_b3_b_122 ), .B (n_8101), .Y (n_8090));
INVX1 g42697(.A (n_444), .Y (n_614));
INVX1 g42690(.A (u9_mem_b2_b_102 ), .Y (n_6635));
INVX2 g35148(.A (n_7402), .Y (n_9055));
INVX1 g35149(.A (n_7402), .Y (n_9036));
INVX1 g35144(.A (n_7402), .Y (n_8976));
INVX1 g35145(.A (n_7402), .Y (n_8951));
INVX1 g35142(.A (n_7402), .Y (n_8948));
INVX1 g35143(.A (n_7402), .Y (n_8961));
INVX1 g35140(.A (n_7402), .Y (n_8958));
INVX1 g35141(.A (n_7402), .Y (n_8971));
OAI21X1 g31045(.A0 (n_5310), .A1 (n_10820), .B0 (n_10364), .Y(n_10866));
INVX1 g42471(.A (n_524), .Y (n_3987));
NAND2X1 g34819(.A (u8_mem_b1_b_69 ), .B (n_7976), .Y (n_7615));
NAND2X1 g34818(.A (u8_mem_b2_b_48 ), .B (n_7976), .Y (n_7616));
INVX1 g42474(.A (u11_mem_b0_b_157 ), .Y (n_6344));
INVX1 g42477(.A (u9_mem_b2_b_117 ), .Y (n_385));
NAND2X1 g34813(.A (u7_mem_b3_b_130 ), .B (n_7651), .Y (n_7620));
NAND2X1 g34812(.A (u7_mem_b3_b_129 ), .B (n_7651), .Y (n_7621));
NAND2X1 g34811(.A (u7_mem_b3_b_128 ), .B (n_7651), .Y (n_7622));
NAND2X1 g34810(.A (u7_mem_b3_b_127 ), .B (n_7651), .Y (n_7623));
NAND2X1 g34817(.A (u3_mem_b2_b_45 ), .B (n_8101), .Y (n_7617));
NAND2X1 g34816(.A (u3_mem_b1_b_63 ), .B (n_8141), .Y (n_7618));
NAND2X1 g34815(.A (u3_mem_b3_b_151 ), .B (n_8097), .Y (n_7619));
NOR2X1 g34814(.A (n_1421), .B (n_7651), .Y (n_8218));
AOI21X1 g35498(.A0 (n_1206), .A1 (i4_re), .B0 (n_6712), .Y (n_7142));
XOR2X1 g35499(.A (n_6049), .B (n_4842), .Y (n_6050));
NAND2X1 g36943(.A (n_2529), .B (n_1317), .Y (n_4811));
NOR2X1 g36942(.A (n_7297), .B (n_4676), .Y (n_5384));
NAND2X1 g36941(.A (n_1638), .B (n_1637), .Y (n_4020));
NAND2X1 g36940(.A (n_1645), .B (n_1642), .Y (n_4021));
AOI21X1 g35360(.A0 (n_6972), .A1 (oc0_cfg_964), .B0 (n_7338), .Y(n_7458));
NAND2X1 g39341(.A (u5_mem_b1_b_67 ), .B (n_3236), .Y (n_12034));
INVX1 g42687(.A (u11_mem_b0_b_156 ), .Y (n_6347));
NAND2X1 g34300(.A (u3_mem_b3_b_136 ), .B (n_8101), .Y (n_8095));
NAND2X1 g39342(.A (n_3259), .B (u5_mem_b0_b_98 ), .Y (n_3261));
CLKBUFX3 g45435(.A (n_11802), .Y (n_11804));
INVX2 g45434(.A (n_11802), .Y (n_11797));
AOI21X1 g38577(.A0 (u8_mem_b2_b_47 ), .A1 (n_4491), .B0 (n_2201), .Y(n_4270));
INVX2 g45436(.A (n_692), .Y (n_11802));
NAND2X1 g39343(.A (u5_mem_b2_b_36 ), .B (n_12823), .Y (n_12035));
AOI21X1 g38257(.A0 (u3_mem_b2_b_42 ), .A1 (n_4519), .B0 (n_2014), .Y(n_4384));
AOI21X1 g38570(.A0 (u7_mem_b3_b_147 ), .A1 (n_5145), .B0 (n_2909), .Y(n_4862));
NAND2X1 g39344(.A (n_3259), .B (u5_mem_b0_b_100 ), .Y (n_3260));
NAND2X1 g36601(.A (n_5798), .B (n_6259), .Y (n_5799));
NAND2X1 g39345(.A (u5_mem_b2_b_38 ), .B (n_12823), .Y (n_12031));
OAI21X1 g33409(.A0 (n_3886), .A1 (n_8894), .B0 (n_8118), .Y (n_8467));
NAND2X1 g34368(.A (n_6068), .B (n_7465), .Y (n_8231));
NAND2X1 g34361(.A (n_6687), .B (n_7466), .Y (n_8232));
NAND2X1 g34360(.A (u4_mem_b1_b_78 ), .B (n_7984), .Y (n_8042));
NAND2X1 g34363(.A (u4_mem_b1_b_79 ), .B (n_7984), .Y (n_8039));
OAI21X1 g33402(.A0 (n_5122), .A1 (n_8856), .B0 (n_8172), .Y (n_8474));
NAND2X1 g34365(.A (u4_mem_b1_b_81 ), .B (n_7984), .Y (n_8036));
OAI21X1 g33404(.A0 (n_4492), .A1 (n_8868), .B0 (n_8171), .Y (n_8472));
NAND2X1 g34367(.A (u4_mem_b1_b_83 ), .B (n_7984), .Y (n_8034));
OAI21X1 g33406(.A0 (n_4493), .A1 (n_8933), .B0 (n_8072), .Y (n_8470));
NAND2X1 g39346(.A (u5_mem_b2_b_35 ), .B (n_12823), .Y (n_2322));
INVX1 g35461(.A (n_7441), .Y (n_863));
AOI21X1 g38468(.A0 (u8_mem_b2_b_55 ), .A1 (n_4499), .B0 (n_1871), .Y(n_4321));
AOI21X1 g38466(.A0 (u6_mem_b2_b_37 ), .A1 (n_4544), .B0 (n_2178), .Y(n_4322));
AOI21X1 g38467(.A0 (u3_mem_b3_b_129 ), .A1 (n_5133), .B0 (n_3329), .Y(n_4908));
AOI21X1 g38464(.A0 (u3_mem_b3_b_139 ), .A1 (n_5138), .B0 (n_2902), .Y(n_4910));
AOI21X1 g38465(.A0 (u7_mem_b3_b_123 ), .A1 (n_5145), .B0 (n_3364), .Y(n_4909));
AOI21X1 g38462(.A0 (u3_mem_b2_b_33 ), .A1 (n_4519), .B0 (n_2029), .Y(n_4324));
AOI21X1 g38463(.A0 (u6_mem_b2_b_30 ), .A1 (n_4504), .B0 (n_1974), .Y(n_4323));
AOI21X1 g38460(.A0 (u8_mem_b3_b_152 ), .A1 (n_3879), .B0 (n_1466), .Y(n_3850));
AOI21X1 g38461(.A0 (u7_mem_b1_b_85 ), .A1 (n_5069), .B0 (n_2711), .Y(n_4911));
NAND2X1 g39347(.A (u5_mem_b1_b_66 ), .B (n_3257), .Y (n_3258));
AOI21X1 g38156(.A0 (u4_mem_b2_b_29 ), .A1 (n_4439), .B0 (n_1827), .Y(n_4429));
AOI21X1 g38253(.A0 (u8_mem_b1_b_80 ), .A1 (n_4387), .B0 (n_2073), .Y(n_4386));
MX2X1 g34033(.A (u5_mem_b0_b_117 ), .B (n_3656), .S0 (n_7496), .Y(n_8792));
AOI21X1 g38208(.A0 (u4_mem_b3_b_146 ), .A1 (n_5102), .B0 (n_3292), .Y(n_5085));
AOI21X1 g38209(.A0 (u6_mem_b2_b_33 ), .A1 (n_4504), .B0 (n_2212), .Y(n_4401));
NAND2X1 g38840(.A (u5_mem_b3_b ), .B (n_1543), .Y (n_1324));
AOI21X1 g38202(.A0 (u4_mem_b3_b_141 ), .A1 (n_5106), .B0 (n_3511), .Y(n_5090));
AOI21X1 g38203(.A0 (u4_mem_b3_b_142 ), .A1 (n_5106), .B0 (n_3295), .Y(n_5089));
AOI21X1 g38200(.A0 (u4_mem_b3_b_140 ), .A1 (n_5106), .B0 (n_3487), .Y(n_5092));
AOI21X1 g38201(.A0 (u4_mem_b3_b_122 ), .A1 (n_5102), .B0 (n_2941), .Y(n_5091));
AOI21X1 g38206(.A0 (u4_mem_b3_b_144 ), .A1 (n_5102), .B0 (n_3293), .Y(n_5087));
AOI21X1 g38207(.A0 (u4_mem_b3_b_145 ), .A1 (n_5102), .B0 (n_3185), .Y(n_5086));
AOI21X1 g38204(.A0 (u4_mem_b3_b_143 ), .A1 (n_5102), .B0 (n_2951), .Y(n_5088));
NAND2X1 g32756(.A (n_103), .B (n_9943), .Y (n_11677));
OR2X1 g32757(.A (n_9512), .B (n_9480), .Y (n_9640));
NAND2X1 g32754(.A (n_191), .B (n_10583), .Y (n_11640));
NAND2X1 g32755(.A (n_183), .B (n_10583), .Y (n_11642));
NAND2X1 g32752(.A (n_359), .B (n_10583), .Y (n_11993));
NAND2X1 g32753(.A (n_372), .B (n_10583), .Y (n_11638));
AOI21X1 g32750(.A0 (n_6245), .A1 (n_6251), .B0 (n_9873), .Y(n_10573));
NAND2X1 g32751(.A (n_322), .B (n_10583), .Y (n_11636));
OR2X1 g32758(.A (n_9511), .B (n_9479), .Y (n_9639));
OR2X1 g32759(.A (n_9510), .B (n_9478), .Y (n_9638));
XOR2X1 g37413(.A (u2_bit_clk_r1), .B (u2_bit_clk_r), .Y (n_2589));
NOR2X1 g39024(.A (n_3332), .B (n_2744), .Y (n_3505));
AOI21X1 g37265(.A0 (n_5492), .A1 (n_6649), .B0 (n_4649), .Y (n_5493));
NAND2X1 g38944(.A (u8_mem_b3_b_137 ), .B (n_2468), .Y (n_2399));
NAND2X1 g38947(.A (u3_mem_b3_b_125 ), .B (n_1517), .Y (n_1518));
NAND2X1 g39027(.A (u6_mem_b1_b_68 ), .B (n_12169), .Y (n_4246));
NAND2X1 g38941(.A (u5_mem_b3_b_148 ), .B (n_3543), .Y (n_3528));
NAND2X1 g38940(.A (u4_mem_b3_b_129 ), .B (n_3546), .Y (n_3529));
NAND2X1 g36437(.A (n_6254), .B (n_12531), .Y (n_6255));
NAND2X1 g36433(.A (n_6800), .B (n_12531), .Y (n_6801));
NAND2X1 g36432(.A (n_6803), .B (n_12357), .Y (n_6804));
NAND2X1 g36431(.A (n_6805), .B (n_12357), .Y (n_6806));
NAND2X1 g36430(.A (n_6807), .B (n_12531), .Y (n_6808));
NAND2X1 g36439(.A (n_6252), .B (n_12531), .Y (n_6253));
NAND2X1 g36438(.A (n_6797), .B (u4_rp_b0_b ), .Y (n_11540));
MX2X1 g36129(.A (n_6411), .B (n_6570), .S0 (n_832), .Y (n_6412));
MX2X1 g36128(.A (n_6453), .B (n_6413), .S0 (n_6649), .Y (n_6414));
NOR2X1 g39026(.A (n_3453), .B (n_2741), .Y (n_3501));
NAND2X1 g36641(.A (n_5270), .B (n_3975), .Y (n_5787));
MX2X1 g36121(.A (n_6478), .B (n_6428), .S0 (n_6649), .Y (n_6429));
MX2X1 g36120(.A (n_5969), .B (n_5983), .S0 (n_5312), .Y (n_5970));
MX2X1 g36123(.A (n_6510), .B (n_6424), .S0 (n_6649), .Y (n_6425));
MX2X1 g36122(.A (n_6473), .B (n_6426), .S0 (n_6649), .Y (n_6427));
MX2X1 g36125(.A (n_6459), .B (n_6419), .S0 (n_6649), .Y (n_6420));
MX2X1 g36124(.A (n_6465), .B (n_6421), .S0 (n_6649), .Y (n_6422));
MX2X1 g36127(.A (n_6415), .B (n_6576), .S0 (n_5407), .Y (n_6416));
MX2X1 g36126(.A (n_6444), .B (n_6417), .S0 (n_6649), .Y (n_6418));
INVX8 g41664(.A (n_1108), .Y (n_3622));
NAND2X1 g36391(.A (n_6176), .B (n_6316), .Y (n_6283));
NAND2X1 g36644(.A (n_5266), .B (n_3974), .Y (n_5785));
NAND2X1 g36645(.A (n_5265), .B (n_2582), .Y (n_5784));
OAI21X1 g36646(.A0 (n_4595), .A1 (n_5213), .B0 (n_6131), .Y (n_6123));
NAND2X1 g39528(.A (n_2330), .B (u7_mem_b0_b_101 ), .Y (n_2291));
NAND2X1 g36647(.A (n_5263), .B (n_3971), .Y (n_5783));
NOR2X1 g39529(.A (n_4996), .B (n_2794), .Y (n_3114));
NOR2X1 g39838(.A (n_3453), .B (n_2755), .Y (n_2930));
NAND2X1 g39839(.A (n_2344), .B (in_slt_430), .Y (n_2241));
AOI22X1 g35507(.A0 (n_5630), .A1 (u2_to_cnt_b5_b ), .B0 (n_5629), .B1(n_4853), .Y (n_6046));
NAND2X1 g39524(.A (u3_mem_b2_b_45 ), .B (n_12619), .Y (n_3119));
AOI21X1 g30878(.A0 (n_11613), .A1 (n_11614), .B0 (n_11033), .Y(n_11040));
AOI21X1 g38512(.A0 (u8_mem_b3_b_135 ), .A1 (n_3879), .B0 (n_1464), .Y(n_3845));
NAND2X1 g39835(.A (n_2491), .B (u7_mem_b0_b_95 ), .Y (n_2473));
NOR2X1 g39832(.A (n_3117), .B (n_2755), .Y (n_2934));
NAND2X1 g39521(.A (u3_mem_b2_b_58 ), .B (n_3330), .Y (n_3122));
NAND2X1 g36446(.A (n_5874), .B (n_6091), .Y (n_5888));
NOR2X1 g39522(.A (n_3332), .B (n_2818), .Y (n_3121));
NAND2X1 g39831(.A (u5_mem_b2_b_41 ), .B (n_12823), .Y (n_12856));
NOR2X1 g39304(.A (n_5102), .B (n_2684), .Y (n_3293));
XOR2X1 g35486(.A (u11_wp_b3_b ), .B (n_1233), .Y (n_4102));
AOI22X1 g35505(.A0 (n_5630), .A1 (n_1819), .B0 (n_5629), .B1(n_1820), .Y (n_5445));
NAND2X1 g36447(.A (n_2565), .B (n_4836), .Y (n_6059));
NAND2X1 g39307(.A (n_12369), .B (u6_mem_b0_b_113 ), .Y (n_3290));
NAND2X1 g39300(.A (u4_mem_b2_b_49 ), .B (n_12091), .Y (n_3297));
NOR2X1 g39301(.A (n_3332), .B (n_2786), .Y (n_3296));
NAND2X1 g39650(.A (u4_mem_b1_b_68 ), .B (n_12252), .Y (n_11663));
AOI21X1 g35480(.A0 (i3_re), .A1 (u9_rp_b2_b ), .B0 (n_6713), .Y(n_7147));
AOI21X1 g30871(.A0 (n_10601), .A1 (n_10504), .B0 (n_5839), .Y(n_11051));
AOI21X1 g30870(.A0 (n_11919), .A1 (n_11724), .B0 (n_5839), .Y(n_11052));
AOI21X1 g30873(.A0 (n_12453), .A1 (n_12672), .B0 (n_5839), .Y(n_11047));
AOI21X1 g30872(.A0 (n_10599), .A1 (n_12690), .B0 (n_5839), .Y(n_11049));
AOI21X1 g30875(.A0 (n_10595), .A1 (n_10496), .B0 (n_11043), .Y(n_11044));
AOI21X1 g30874(.A0 (n_12464), .A1 (n_11748), .B0 (n_11043), .Y(n_11045));
AOI21X1 g30877(.A0 (n_10592), .A1 (n_10493), .B0 (n_5839), .Y(n_11041));
AOI21X1 g30876(.A0 (n_11633), .A1 (n_11634), .B0 (n_11030), .Y(n_11042));
AOI21X1 g30879(.A0 (n_11615), .A1 (n_11616), .B0 (n_12585), .Y(n_11039));
NOR2X1 g35809(.A (n_980), .B (n_6752), .Y (n_6739));
NAND2X1 g39527(.A (u4_mem_b1_b_85 ), .B (n_12270), .Y (n_4177));
NOR2X1 g39520(.A (n_4996), .B (n_2767), .Y (n_3123));
NAND2X1 g39833(.A (u7_mem_b1_b_70 ), .B (n_4130), .Y (n_4114));
NAND2X1 g39830(.A (u7_mem_b2_b_48 ), .B (n_12654), .Y (n_3553));
NAND2X1 g39523(.A (u7_mem_b2_b_40 ), .B (n_12645), .Y (n_3120));
INVX1 g42314(.A (u11_mem_b1_b_131 ), .Y (n_6511));
INVX1 g42316(.A (n_4736), .Y (n_936));
AOI21X1 g34178(.A0 (n_1417), .A1 (n_7758), .B0 (n_8221), .Y (n_9361));
AOI21X1 g34179(.A0 (n_1421), .A1 (n_7651), .B0 (n_8218), .Y (n_9360));
AOI21X1 g38113(.A0 (u4_mem_b1_b_73 ), .A1 (n_4471), .B0 (n_1961), .Y(n_4467));
AOI21X1 g34174(.A0 (u8_wp_b0_b ), .A1 (n_7976), .B0 (n_8248), .Y(n_9365));
AOI21X1 g34175(.A0 (n_1419), .A1 (n_7984), .B0 (n_8227), .Y (n_9364));
AOI21X1 g34176(.A0 (n_798), .A1 (n_7870), .B0 (n_8224), .Y (n_9363));
AOI21X1 g34177(.A0 (n_1424), .A1 (n_8141), .B0 (n_8241), .Y (n_9362));
MX2X1 g34170(.A (u3_mem_b0_b_96 ), .B (n_3574), .S0 (n_8700), .Y(n_9366));
MX2X1 g34171(.A (u3_mem_b0_b_97 ), .B (n_3654), .S0 (n_7423), .Y(n_8249));
MX2X1 g34172(.A (u3_mem_b0_b_98 ), .B (n_3572), .S0 (n_8700), .Y(n_8681));
MX2X1 g34173(.A (u3_mem_b0_b_99 ), .B (n_3751), .S0 (n_8700), .Y(n_8680));
NAND2X1 g39658(.A (u6_mem_b1_b_87 ), .B (n_4253), .Y (n_4150));
NOR2X1 g39659(.A (n_3117), .B (n_2829), .Y (n_2739));
AOI21X1 g38289(.A0 (u5_mem_b1_b_71 ), .A1 (n_5048), .B0 (n_2816), .Y(n_5023));
AOI21X1 g38114(.A0 (u7_mem_b2_b_46 ), .A1 (n_4509), .B0 (n_2000), .Y(n_4466));
NAND2X1 g36933(.A (n_2532), .B (n_1237), .Y (n_4813));
NAND2X1 g39788(.A (n_12825), .B (u3_mem_b0_b_112 ), .Y (n_2957));
NAND2X1 g39789(.A (n_2330), .B (u7_mem_b0_b_104 ), .Y (n_2489));
NAND2X1 g36931(.A (n_1662), .B (n_1661), .Y (n_4027));
NAND2X1 g38899(.A (u6_mem_b3_b_123 ), .B (n_12622), .Y (n_2414));
NAND2X1 g39780(.A (n_2325), .B (in_slt_448), .Y (n_2248));
NAND2X1 g39781(.A (u7_mem_b1_b_71 ), .B (n_4130), .Y (n_4127));
NOR2X1 g39782(.A (n_5102), .B (n_2765), .Y (n_2962));
NOR2X1 g39783(.A (n_3089), .B (n_2729), .Y (n_2961));
NAND2X1 g39784(.A (u7_mem_b2_b_53 ), .B (n_12650), .Y (n_4126));
NAND2X1 g39785(.A (n_3252), .B (u7_mem_b0_b_103 ), .Y (n_2959));
NAND2X1 g39786(.A (n_2491), .B (u7_mem_b0_b_108 ), .Y (n_2247));
NOR2X1 g39787(.A (n_5102), .B (n_2767), .Y (n_2958));
XOR2X1 g35501(.A (n_5618), .B (n_4091), .Y (n_5619));
MX2X1 g36026(.A (n_6602), .B (n_6601), .S0 (n_6594), .Y (n_6603));
NOR2X1 g40923(.A (u11_wp_b1_b ), .B (n_520), .Y (n_932));
NAND2X1 g36938(.A (n_1651), .B (n_1648), .Y (n_4023));
INVX8 g40925(.A (n_1162), .Y (n_5341));
NAND2X1 g39029(.A (u3_mem_b1_b_83 ), .B (n_3316), .Y (n_3499));
OAI21X1 g31043(.A0 (n_5311), .A1 (n_10820), .B0 (n_10365), .Y(n_10867));
OAI21X1 g31042(.A0 (n_5322), .A1 (n_10820), .B0 (n_10366), .Y(n_10868));
NAND3X1 g31737(.A (n_6816), .B (n_10518), .C (n_1873), .Y (n_11109));
NAND2X1 g39028(.A (u6_mem_b1_b_88 ), .B (n_4253), .Y (n_4244));
OAI21X1 g31040(.A0 (n_5316), .A1 (n_10820), .B0 (n_10369), .Y(n_10872));
AND2X1 g31731(.A (n_5626), .B (ac97_rst_force), .Y (n_9493));
NAND2X1 g31730(.A (n_5522), .B (n_10385), .Y (n_10345));
INVX4 g32929(.A (n_9721), .Y (n_9820));
AOI21X1 g31733(.A0 (n_2369), .A1 (n_4829), .B0 (n_11894), .Y(n_9974));
OAI21X1 g31044(.A0 (n_5408), .A1 (n_10450), .B0 (n_9988), .Y(n_10676));
NOR2X1 g40229(.A (n_2782), .B (n_2067), .Y (n_2022));
NOR2X1 g40228(.A (n_2154), .B (n_2801), .Y (n_2023));
NOR2X1 g40227(.A (n_2477), .B (n_3008), .Y (n_2024));
NOR2X1 g40226(.A (n_2705), .B (n_2735), .Y (n_2706));
AOI22X1 g37988(.A0 (n_2502), .A1 (n_6845), .B0 (n_6937), .B1(n_1859), .Y (n_2498));
NAND2X1 g40224(.A (n_4507), .B (n_4439), .Y (n_1450));
NOR2X1 g40223(.A (n_2071), .B (n_2686), .Y (n_2027));
NOR2X1 g40222(.A (n_2829), .B (n_933), .Y (n_2028));
NOR2X1 g40221(.A (n_2071), .B (n_2744), .Y (n_2029));
NOR2X1 g40220(.A (n_1147), .B (n_2707), .Y (n_2709));
NAND2X1 g39579(.A (n_12369), .B (u6_mem_b0_b_114 ), .Y (n_3086));
NAND2X1 g32696(.A (n_212), .B (n_10617), .Y (n_10623));
NAND2X1 g32695(.A (n_181), .B (n_10617), .Y (n_10625));
NAND2X1 g32694(.A (n_167), .B (n_10617), .Y (n_10626));
NAND2X1 g32693(.A (n_10617), .B (n_1481), .Y (n_11104));
NAND2X1 g32692(.A (n_243), .B (n_9943), .Y (n_12001));
NAND2X1 g32691(.A (n_332), .B (n_9943), .Y (n_12011));
NAND2X1 g32690(.A (n_10787), .B (n_991), .Y (n_10953));
OAI21X1 g32699(.A0 (n_5594), .A1 (n_7529), .B0 (n_7528), .Y (n_7530));
NAND2X1 g32698(.A (n_76), .B (n_10617), .Y (n_10622));
NOR2X1 g40322(.A (n_2470), .B (n_2702), .Y (n_1962));
NOR2X1 g40323(.A (n_2470), .B (n_2755), .Y (n_1961));
NOR2X1 g40320(.A (n_2770), .B (n_2790), .Y (n_2669));
NOR2X1 g40321(.A (n_2696), .B (n_2702), .Y (n_2668));
NOR2X1 g40326(.A (n_2759), .B (n_2702), .Y (n_2665));
NOR2X1 g40327(.A (n_2689), .B (n_2732), .Y (n_2664));
NOR2X1 g40324(.A (n_1082), .B (n_2792), .Y (n_2667));
OAI21X1 g45941(.A0 (n_12683), .A1 (n_12686), .B0 (n_12689), .Y(n_12690));
INVX1 g45940(.A (n_12678), .Y (n_12682));
NOR2X1 g40328(.A (n_2741), .B (n_2045), .Y (n_1960));
NOR2X1 g40329(.A (n_2742), .B (n_2790), .Y (n_2663));
NAND2X1 g45945(.A (n_12115), .B (n_12116), .Y (n_12685));
NAND2X1 g45944(.A (n_12664), .B (n_12111), .Y (n_12684));
NAND2X1 g39330(.A (n_3259), .B (u5_mem_b0_b ), .Y (n_3270));
INVX4 g45946(.A (n_12688), .Y (n_12689));
AOI21X1 g38071(.A0 (u3_mem_b3_b_126 ), .A1 (n_5133), .B0 (n_2880), .Y(n_5125));
AOI21X1 g38070(.A0 (u8_mem_b2_b_43 ), .A1 (n_4491), .B0 (n_1884), .Y(n_4495));
AOI21X1 g38073(.A0 (u8_mem_b2_b_42 ), .A1 (n_4499), .B0 (n_1993), .Y(n_4494));
AOI21X1 g38075(.A0 (u3_mem_b3_b_128 ), .A1 (n_5138), .B0 (n_3370), .Y(n_5124));
AOI21X1 g38074(.A0 (u8_mem_b2_b_36 ), .A1 (n_4499), .B0 (n_2183), .Y(n_4493));
AOI21X1 g38077(.A0 (u3_mem_b3_b_148 ), .A1 (n_5133), .B0 (n_3865), .Y(n_5123));
AOI21X1 g38076(.A0 (u8_mem_b2_b_35 ), .A1 (n_4491), .B0 (n_2160), .Y(n_4492));
AOI21X1 g38079(.A0 (u8_mem_b2_b_34 ), .A1 (n_4499), .B0 (n_2174), .Y(n_4490));
AOI21X1 g38078(.A0 (u3_mem_b1_b_88 ), .A1 (n_5148), .B0 (n_2803), .Y(n_5122));
AOI21X1 g38332(.A0 (u5_mem_b2_b_34 ), .A1 (n_4378), .B0 (n_2013), .Y(n_4354));
AOI21X1 g38333(.A0 (u5_mem_b2_b_35 ), .A1 (n_4370), .B0 (n_2015), .Y(n_4353));
AOI21X1 g38330(.A0 (u7_mem_b1_b_87 ), .A1 (n_5069), .B0 (n_2740), .Y(n_5005));
AOI21X1 g38331(.A0 (u6_mem_b1_b_81 ), .A1 (n_5019), .B0 (n_2797), .Y(n_5004));
AOI21X1 g38336(.A0 (u5_mem_b2_b_37 ), .A1 (n_4370), .B0 (n_1980), .Y(n_4351));
MX2X1 g38625(.A (u4_mem_b0_b_114 ), .B (wb_din_684), .S0 (n_3765), .Y(n_3770));
INVX1 g37106(.A (n_6155), .Y (n_5672));
NAND2X1 g34325(.A (u3_mem_b3_b_129 ), .B (n_8141), .Y (n_8073));
NAND4X1 g37107(.A (n_12036), .B (n_1493), .C (n_12037), .D (n_2399),.Y (n_6155));
NOR2X1 g40156(.A (n_2081), .B (n_2763), .Y (n_2082));
MX2X1 g38695(.A (u6_mem_b0_b_99 ), .B (wb_din_669), .S0 (n_3632), .Y(n_3658));
MX2X1 g38694(.A (u6_mem_b0_b_98 ), .B (wb_din_668), .S0 (n_813), .Y(n_3660));
MX2X1 g38697(.A (u3_mem_b0_b_97 ), .B (wb_din_667), .S0 (n_3807), .Y(n_3654));
MX2X1 g38696(.A (u5_mem_b0_b_117 ), .B (wb_din_687), .S0 (n_3720), .Y(n_3656));
MX2X1 g38691(.A (u6_mem_b0_b_121 ), .B (wb_din_691), .S0 (n_3632), .Y(n_3666));
MX2X1 g38690(.A (u6_mem_b0_b_120 ), .B (wb_din_690), .S0 (n_3632), .Y(n_3667));
MX2X1 g38693(.A (u6_mem_b0_b_97 ), .B (wb_din_667), .S0 (n_813), .Y(n_3663));
MX2X1 g38692(.A (u6_mem_b0_b_95 ), .B (wb_din_665), .S0 (n_3632), .Y(n_3664));
MX2X1 g38699(.A (u8_mem_b0_b_117 ), .B (wb_din_687), .S0 (n_3826), .Y(n_3651));
MX2X1 g38698(.A (u6_mem_b0_b_96 ), .B (wb_din_666), .S0 (n_3632), .Y(n_3652));
NAND2X1 g41321(.A (n_5225), .B (wb_addr_i_b4_b), .Y (n_3431));
OR2X1 g41320(.A (n_11563), .B (n_1308), .Y (n_1309));
INVX1 g41325(.A (n_844), .Y (n_1136));
OR2X1 g41326(.A (n_410), .B (n_11578), .Y (n_844));
NAND2X1 g39285(.A (n_3316), .B (u3_mem_b1_b_72 ), .Y (n_3317));
NAND2X1 g38888(.A (u6_mem_b3_b_128 ), .B (n_2419), .Y (n_2426));
NAND2X1 g36334(.A (n_5713), .B (n_6318), .Y (n_6314));
NAND2X1 g36335(.A (n_5561), .B (n_6318), .Y (n_5932));
NAND2X1 g36336(.A (n_5863), .B (n_6318), .Y (n_5931));
NAND2X1 g36330(.A (n_5886), .B (n_6318), .Y (n_5936));
NAND2X1 g36331(.A (n_5884), .B (n_6318), .Y (n_5935));
NAND2X1 g36332(.A (n_5882), .B (n_6318), .Y (n_5934));
NAND2X1 g36333(.A (n_5879), .B (n_6318), .Y (n_5933));
NAND2X1 g40810(.A (n_37), .B (u26_cnt_b2_b ), .Y (n_713));
NOR2X1 g40811(.A (n_2567), .B (u8_rp_b3_b ), .Y (n_639));
MX2X1 g31319(.A (n_6358), .B (n_6357), .S0 (n_10537), .Y (n_10430));
NAND2X1 g31649(.A (n_5369), .B (n_10019), .Y (n_9997));
OR2X1 g31648(.A (n_10329), .B (n_765), .Y (n_9998));
NAND2X1 g40816(.A (n_53), .B (u9_rp_b0_b ), .Y (n_877));
INVX1 g40817(.A (n_806), .Y (n_6141));
MX2X1 g31313(.A (n_5660), .B (n_1600), .S0 (n_10513), .Y (n_10436));
MX2X1 g31312(.A (n_5650), .B (n_1605), .S0 (n_10537), .Y (n_10437));
MX2X1 g31311(.A (n_5472), .B (n_1244), .S0 (n_9724), .Y (n_10438));
MX2X1 g31310(.A (n_5651), .B (n_1610), .S0 (n_10537), .Y (n_10439));
MX2X1 g31317(.A (n_5649), .B (n_1242), .S0 (n_10137), .Y (n_10129));
MX2X1 g31316(.A (n_5658), .B (n_1592), .S0 (n_10537), .Y (n_10432));
MX2X1 g31315(.A (n_5644), .B (n_1596), .S0 (n_10513), .Y (n_10433));
MX2X1 g31314(.A (n_5662), .B (n_2557), .S0 (n_9724), .Y (n_10435));
XOR2X1 g37422(.A (n_6841), .B (n_754), .Y (n_1265));
XOR2X1 g37421(.A (n_7048), .B (n_762), .Y (n_1267));
XOR2X1 g37420(.A (n_657), .B (n_771), .Y (n_1788));
NOR2X1 g41499(.A (u11_wp_b1_b ), .B (n_853), .Y (n_1072));
NAND2X1 g39287(.A (u3_mem_b2_b_50 ), .B (n_3330), .Y (n_3315));
INVX8 g41496(.A (n_1854), .Y (n_6359));
INVX2 g41494(.A (n_1072), .Y (n_1854));
NAND2X1 g35831(.A (n_1815), .B (n_5248), .Y (n_5249));
INVX1 g42107(.A (u8_rp_b1_b ), .Y (n_244));
NAND2X1 g36590(.A (n_5807), .B (n_6259), .Y (n_5808));
NAND2X1 g36591(.A (n_6165), .B (n_634), .Y (n_6166));
NAND2X1 g36592(.A (n_6163), .B (n_12115), .Y (n_6164));
NAND2X1 g36593(.A (n_5805), .B (n_6259), .Y (n_5806));
NAND2X1 g36594(.A (n_6161), .B (n_12115), .Y (n_6162));
NAND2X1 g36595(.A (n_6159), .B (n_6259), .Y (n_6160));
NAND2X1 g36596(.A (n_5803), .B (n_1038), .Y (n_5804));
NAND2X1 g36597(.A (n_6157), .B (n_12115), .Y (n_6158));
NAND2X1 g36598(.A (n_6155), .B (n_6152), .Y (n_6156));
NAND2X1 g36599(.A (n_5800), .B (n_6259), .Y (n_5801));
INVX1 g36983(.A (n_6786), .Y (n_6074));
INVX1 g42678(.A (u9_mem_b0_b_150 ), .Y (n_6862));
INVX1 g42676(.A (u10_mem_b2_b_113 ), .Y (n_379));
INVX1 g42674(.A (oc2_cfg_987), .Y (n_503));
OAI21X1 g30998(.A0 (n_5370), .A1 (n_10747), .B0 (n_9997), .Y(n_10705));
OAI21X1 g30999(.A0 (n_5368), .A1 (n_10738), .B0 (n_10018), .Y(n_10704));
OAI21X1 g30992(.A0 (n_5295), .A1 (n_10747), .B0 (n_10027), .Y(n_10711));
OAI21X1 g30993(.A0 (n_5375), .A1 (n_10747), .B0 (n_10026), .Y(n_10710));
OAI21X1 g30990(.A0 (n_6090), .A1 (n_10738), .B0 (n_10029), .Y(n_10713));
OAI21X1 g30991(.A0 (n_6088), .A1 (n_10747), .B0 (n_10028), .Y(n_10712));
OAI21X1 g30996(.A0 (n_5334), .A1 (n_10747), .B0 (n_10022), .Y(n_10707));
OAI21X1 g30997(.A0 (n_5303), .A1 (n_10747), .B0 (n_10020), .Y(n_10706));
OAI21X1 g30994(.A0 (n_5344), .A1 (n_10019), .B0 (n_10025), .Y(n_10709));
OAI21X1 g30995(.A0 (n_5373), .A1 (n_10747), .B0 (n_10023), .Y(n_10708));
INVX1 g45378(.A (n_11597), .Y (n_11600));
NOR2X1 g39282(.A (n_3453), .B (n_2748), .Y (n_3321));
INVX1 g42411(.A (u11_mem_b0_b_160 ), .Y (n_6370));
INVX1 g42416(.A (u11_mem_b2_b_105 ), .Y (n_129));
INVX1 g42414(.A (u9_mem_b1_b_137 ), .Y (n_1748));
INVX1 g42415(.A (u11_mem_b0_b_170 ), .Y (n_1628));
AOI21X1 g35344(.A0 (i4_dout_597), .A1 (n_7468), .B0 (n_7346), .Y(n_7469));
AOI21X1 g35345(.A0 (i4_dout_598), .A1 (n_7468), .B0 (n_7345), .Y(n_7467));
AOI21X1 g35346(.A0 (i4_dout_599), .A1 (n_7468), .B0 (n_7344), .Y(n_7466));
AOI21X1 g35347(.A0 (i4_dout_600), .A1 (n_7468), .B0 (n_7343), .Y(n_7465));
AOI21X1 g35340(.A0 (i4_dout_605), .A1 (n_7468), .B0 (n_7351), .Y(n_7473));
AOI21X1 g35341(.A0 (i4_dout_606), .A1 (n_7468), .B0 (n_7350), .Y(n_7472));
AOI21X1 g35342(.A0 (i4_dout_609), .A1 (n_7468), .B0 (n_7354), .Y(n_7471));
AOI21X1 g35343(.A0 (i4_dout_596), .A1 (n_7468), .B0 (n_7347), .Y(n_7470));
NAND2X1 g39319(.A (n_4560), .B (in_slt_453), .Y (n_5280));
INVX1 g39318(.A (n_5280), .Y (n_4202));
AOI21X1 g35348(.A0 (i4_dout_601), .A1 (n_7468), .B0 (n_7342), .Y(n_7464));
AOI21X1 g35349(.A0 (i4_dout_602), .A1 (n_7468), .B0 (n_7341), .Y(n_7463));
NAND4X1 g36921(.A (n_11439), .B (n_3193), .C (n_11440), .D (n_2438),.Y (n_5865));
NAND2X1 g36923(.A (n_1668), .B (n_1667), .Y (n_4030));
NAND2X1 g36922(.A (n_2543), .B (n_1252), .Y (n_4814));
NAND2X1 g36927(.A (n_1666), .B (n_1891), .Y (n_4029));
NAND4X1 g36926(.A (n_12809), .B (n_12810), .C (n_2560), .D (n_1337),.Y (n_5707));
NOR2X1 g36929(.A (n_1025), .B (n_2513), .Y (n_2606));
NAND4X1 g36928(.A (n_3526), .B (n_3186), .C (n_3288), .D (n_1791), .Y(n_5557));
NAND2X1 g38880(.A (u4_mem_b3_b_132 ), .B (n_12744), .Y (n_11655));
NOR2X1 g34699(.A (n_1417), .B (n_7758), .Y (n_8221));
NAND2X1 g34698(.A (u8_mem_b3_b_152 ), .B (n_7976), .Y (n_7727));
NOR2X1 g37585(.A (n_5298), .B (n_6649), .Y (n_4636));
NAND2X1 g34691(.A (u6_mem_b3_b_125 ), .B (n_7758), .Y (n_7733));
NAND2X1 g34690(.A (u6_mem_b3_b_124 ), .B (n_7758), .Y (n_7734));
NOR2X1 g34693(.A (o7_status_992), .B (n_422), .Y (n_9546));
NAND2X1 g34692(.A (u6_mem_b3_b_126 ), .B (n_7758), .Y (n_7732));
NAND2X1 g34695(.A (u6_mem_b3_b_128 ), .B (n_7758), .Y (n_7730));
NAND2X1 g34694(.A (u6_mem_b3_b_127 ), .B (n_7758), .Y (n_7731));
NAND2X1 g34697(.A (u6_mem_b3_b_130 ), .B (n_7758), .Y (n_7728));
NAND2X1 g34696(.A (u6_mem_b3_b_129 ), .B (n_7758), .Y (n_7729));
AND2X1 g37587(.A (n_2412), .B (n_3944), .Y (n_3945));
NOR2X1 g37583(.A (n_5335), .B (n_6649), .Y (n_4638));
OAI21X1 g33423(.A0 (n_3869), .A1 (n_8894), .B0 (n_8047), .Y (n_8446));
OAI21X1 g33422(.A0 (n_5151), .A1 (n_8097), .B0 (n_7818), .Y (n_8447));
OAI21X1 g33421(.A0 (n_3871), .A1 (n_8449), .B0 (n_8156), .Y (n_8448));
OAI21X1 g33420(.A0 (n_3843), .A1 (n_8449), .B0 (n_8157), .Y (n_8450));
NAND2X1 g34431(.A (u4_mem_b3_b_131 ), .B (n_7984), .Y (n_7985));
OAI21X1 g33426(.A0 (n_3874), .A1 (n_8453), .B0 (n_8152), .Y (n_8442));
NAND2X1 g34433(.A (u8_mem_b1_b ), .B (n_7976), .Y (n_7982));
NAND2X1 g34432(.A (u4_mem_b3_b_132 ), .B (n_7984), .Y (n_7983));
OAI21X1 g33429(.A0 (n_3880), .A1 (n_8438), .B0 (n_8150), .Y (n_8437));
OAI21X1 g33428(.A0 (n_3878), .A1 (n_8438), .B0 (n_8151), .Y (n_8439));
NAND2X1 g34439(.A (u4_mem_b3_b_137 ), .B (n_7984), .Y (n_7975));
NAND2X1 g34438(.A (u8_mem_b2_b_56 ), .B (n_7976), .Y (n_7977));
NAND2X1 g39288(.A (u5_mem_b1_b_63 ), .B (n_3236), .Y (n_12800));
NAND2X1 g36506(.A (n_5829), .B (n_6816), .Y (n_5846));
AOI21X1 g38448(.A0 (u6_mem_b3_b_123 ), .A1 (n_5059), .B0 (n_3285), .Y(n_4919));
AOI21X1 g38449(.A0 (u8_mem_b2_b_54 ), .A1 (n_4491), .B0 (n_1986), .Y(n_4326));
AOI21X1 g38198(.A0 (u4_mem_b3_b_139 ), .A1 (n_5102), .B0 (n_3299), .Y(n_5094));
AOI21X1 g38199(.A0 (u3_mem_b3_b_143 ), .A1 (n_5138), .B0 (n_2954), .Y(n_5093));
AOI21X1 g38440(.A0 (u6_mem_b3_b_134 ), .A1 (n_5059), .B0 (n_2946), .Y(n_4925));
AOI21X1 g38193(.A0 (u4_mem_b3_b_136 ), .A1 (n_5106), .B0 (n_3305), .Y(n_5098));
AOI21X1 g38190(.A0 (u6_mem_b3_b_126 ), .A1 (n_5100), .B0 (n_3505), .Y(n_5101));
AOI21X1 g38191(.A0 (u4_mem_b3_b_135 ), .A1 (n_5102), .B0 (n_3844), .Y(n_5099));
AOI21X1 g38445(.A0 (u6_mem_b3_b_140 ), .A1 (n_5059), .B0 (n_3121), .Y(n_4922));
AOI21X1 g38194(.A0 (u6_mem_b1_b_63 ), .A1 (n_5112), .B0 (n_2796), .Y(n_5097));
AOI21X1 g38195(.A0 (u4_mem_b3_b_137 ), .A1 (n_5106), .B0 (n_3434), .Y(n_5096));
INVX1 g42833(.A (u9_mem_b2_b_103 ), .Y (n_6873));
INVX1 g42834(.A (u11_mem_b0_b_155 ), .Y (n_6349));
NAND2X1 g34354(.A (u4_mem_b1_b_73 ), .B (n_7984), .Y (n_8049));
NAND2X1 g34427(.A (u4_mem_b2_b_35 ), .B (n_7984), .Y (n_7989));
NAND2X1 g34424(.A (u4_mem_b2_b_32 ), .B (n_7984), .Y (n_7992));
OAI21X1 g33431(.A0 (n_3881), .A1 (n_8438), .B0 (n_8149), .Y (n_8435));
NOR2X1 g34893(.A (n_7365), .B (n_4800), .Y (n_7512));
NOR2X1 g34892(.A (o9_status), .B (o9_status_1012), .Y (n_7163));
CLKBUFX3 g45429(.A (n_11802), .Y (n_11789));
NOR2X1 g34891(.A (o8_status), .B (o8_status_1002), .Y (n_7164));
OAI21X1 g33699(.A0 (n_4965), .A1 (n_9202), .B0 (n_7840), .Y (n_9198));
NOR2X1 g34890(.A (o7_status), .B (o7_status_992), .Y (n_7165));
NAND3X1 g34897(.A (n_7493), .B (n_2052), .C (n_1481), .Y (n_8673));
NAND2X1 g34724(.A (u7_mem_b1_b_76 ), .B (n_7651), .Y (n_7712));
INVX8 g32772(.A (n_9749), .Y (n_10747));
INVX2 g32774(.A (n_10024), .Y (n_9749));
NAND3X1 g34895(.A (n_7505), .B (n_1972), .C (n_1873), .Y (n_8674));
MX2X1 g38641(.A (u8_mem_b0_b_96 ), .B (wb_din_666), .S0 (n_3826), .Y(n_3750));
OAI21X1 g33438(.A0 (n_3855), .A1 (n_8930), .B0 (n_8140), .Y (n_8426));
NAND3X1 g34894(.A (n_8700), .B (n_2157), .C (n_862), .Y (n_8675));
NOR2X1 g40349(.A (n_2059), .B (n_2729), .Y (n_1945));
OAI21X1 g33439(.A0 (n_3860), .A1 (n_8433), .B0 (n_8139), .Y (n_8425));
NAND2X1 g39598(.A (n_12679), .B (u5_mem_b0_b_114 ), .Y (n_3071));
NOR2X1 g40082(.A (n_2133), .B (n_2804), .Y (n_2152));
AOI21X1 g38225(.A0 (u4_mem_b3_b_126 ), .A1 (n_5106), .B0 (n_3525), .Y(n_5071));
AOI21X1 g38226(.A0 (u7_mem_b1_b_65 ), .A1 (n_5069), .B0 (n_2766), .Y(n_5070));
AOI21X1 g38227(.A0 (u4_mem_b3_b_127 ), .A1 (n_5102), .B0 (n_2962), .Y(n_5068));
AOI21X1 g38220(.A0 (u7_mem_b3_b_138 ), .A1 (n_4961), .B0 (n_3163), .Y(n_5076));
AOI21X1 g38221(.A0 (u4_mem_b3_b_152 ), .A1 (n_5106), .B0 (n_3279), .Y(n_5075));
AOI21X1 g38222(.A0 (u4_mem_b3_b_124 ), .A1 (n_5106), .B0 (n_3280), .Y(n_5074));
AOI21X1 g38223(.A0 (u7_mem_b3_b_143 ), .A1 (n_5145), .B0 (n_3535), .Y(n_5073));
OR2X1 g38998(.A (n_605), .B (n_2368), .Y (n_2371));
NAND2X1 g38999(.A (u8_mem_b3_b_130 ), .B (n_2468), .Y (n_2370));
AOI21X1 g38229(.A0 (u3_mem_b3_b_150 ), .A1 (n_5133), .B0 (n_3463), .Y(n_5066));
MX2X1 g36103(.A (n_6460), .B (n_6459), .S0 (n_5312), .Y (n_6461));
MX2X1 g36102(.A (n_6463), .B (n_6596), .S0 (n_5407), .Y (n_6464));
MX2X1 g36101(.A (n_6466), .B (n_6465), .S0 (n_5409), .Y (n_6467));
MX2X1 g36100(.A (n_6468), .B (n_6599), .S0 (n_5407), .Y (n_6469));
MX2X1 g36107(.A (n_502), .B (n_6586), .S0 (n_6475), .Y (n_6452));
MX2X1 g36106(.A (n_6454), .B (n_6453), .S0 (n_932), .Y (n_6455));
NAND2X1 g36457(.A (n_6241), .B (n_5881), .Y (n_6243));
NAND2X1 g36458(.A (n_5874), .B (n_6141), .Y (n_5875));
MX2X1 g36109(.A (n_6533), .B (n_6450), .S0 (n_6908), .Y (n_6451));
MX2X1 g36108(.A (n_5974), .B (n_6014), .S0 (n_6475), .Y (n_5975));
NOR2X1 g39591(.A (n_4961), .B (n_2729), .Y (n_3076));
NOR2X1 g41289(.A (u13_ints_r_b6_b ), .B (n_540), .Y (n_541));
NAND2X1 g39590(.A (n_12840), .B (u4_mem_b0_b ), .Y (n_11670));
MX2X1 g38628(.A (u4_mem_b0_b_117 ), .B (wb_din_687), .S0 (n_3765), .Y(n_3764));
NAND2X1 g39593(.A (u8_mem_b1_b_90 ), .B (n_12291), .Y (n_3074));
MX2X1 g38629(.A (u4_mem_b0_b_118 ), .B (wb_din_688), .S0 (n_835), .Y(n_3763));
NAND2X1 g40745(.A (n_12281), .B (u8_rp_b1_b ), .Y (n_637));
NAND2X1 g45526(.A (n_6824), .B (n_6805), .Y (n_12131));
INVX2 g41285(.A (n_12535), .Y (n_7214));
NAND2X1 g37856(.A (n_4224), .B (n_3437), .Y (n_12050));
NAND4X1 g37360(.A (n_792), .B (n_549), .C (n_728), .D (n_543), .Y(n_1794));
AOI22X1 g37855(.A0 (n_6434), .A1 (n_1575), .B0 (n_6658), .B1(n_1831), .Y (n_1571));
AOI22X1 g37852(.A0 (n_1756), .A1 (n_6349), .B0 (n_6487), .B1(n_1643), .Y (n_1572));
NAND2X1 g37853(.A (n_2448), .B (n_2955), .Y (n_12049));
NAND2X1 g37850(.A (n_4167), .B (n_3290), .Y (n_12056));
AOI22X1 g37851(.A0 (n_6437), .A1 (n_1575), .B0 (n_6556), .B1(n_1831), .Y (n_1573));
NAND2X1 g38802(.A (u4_mem_b3_b_143 ), .B (n_3556), .Y (n_3557));
NAND2X1 g37858(.A (n_4117), .B (n_1565), .Y (n_5205));
NAND2X1 g37859(.A (n_2440), .B (n_3424), .Y (n_12053));
MX2X1 g33166(.A (wb_din_667), .B (oc0_cfg_970), .S0 (n_8538), .Y(n_8524));
MX2X1 g33167(.A (wb_din_668), .B (n_991), .S0 (n_8538), .Y (n_8523));
MX2X1 g33164(.A (wb_din_665), .B (n_8526), .S0 (n_8538), .Y (n_8527));
MX2X1 g33165(.A (wb_din_666), .B (oc0_cfg_969), .S0 (n_8538), .Y(n_8525));
MX2X1 g33162(.A (wb_din_663), .B (oc0_cfg_966), .S0 (n_8538), .Y(n_8530));
MX2X1 g33163(.A (wb_din_664), .B (n_8528), .S0 (n_8538), .Y (n_8529));
MX2X1 g33160(.A (wb_din_690), .B (oc3_cfg_999), .S0 (n_8538), .Y(n_8534));
MX2X1 g33161(.A (wb_din_691), .B (oc3_cfg_1000), .S0 (n_8538), .Y(n_8532));
NAND2X1 g38804(.A (u8_mem_b3_b_131 ), .B (n_2468), .Y (n_2457));
MX2X1 g33168(.A (wb_din_669), .B (oc1_cfg_974), .S0 (n_8538), .Y(n_8522));
MX2X1 g33169(.A (wb_din), .B (n_1481), .S0 (n_8202), .Y (n_8204));
OAI21X1 g32697(.A0 (n_5595), .A1 (n_7532), .B0 (n_7531), .Y (n_7533));
NAND2X1 g37722(.A (n_2923), .B (n_3159), .Y (n_4601));
INVX1 g42080(.A (u9_mem_b1_b_125 ), .Y (n_6940));
INVX1 g42082(.A (u9_mem_b1_b_141 ), .Y (n_340));
AOI22X1 g37367(.A0 (n_5272), .A1 (u13_intm_r_b11_b ), .B0 (n_5277),.B1 (crac_din_702), .Y (n_5252));
INVX1 g42088(.A (u9_mem_b1_b_126 ), .Y (n_6537));
NAND4X1 g37368(.A (n_732), .B (n_557), .C (n_574), .D (n_725), .Y(n_1793));
INVX1 g45494(.A (n_12079), .Y (n_12077));
AOI21X1 g38575(.A0 (u8_mem_b2_b_53 ), .A1 (n_4491), .B0 (n_2192), .Y(n_4271));
MX2X1 g31108(.A (n_6948), .B (n_6947), .S0 (n_10308), .Y (n_10299));
MX2X1 g31109(.A (n_6877), .B (n_6876), .S0 (n_10308), .Y (n_10298));
MX2X1 g31107(.A (n_6880), .B (n_6879), .S0 (n_10250), .Y (n_10300));
MX2X1 g31104(.A (n_6955), .B (n_6954), .S0 (n_10303), .Y (n_10304));
MX2X1 g31105(.A (n_6950), .B (n_6949), .S0 (n_10250), .Y (n_10302));
MX2X1 g31102(.A (n_6529), .B (n_6528), .S0 (n_10308), .Y (n_10306));
MX2X1 g31103(.A (n_6885), .B (n_6884), .S0 (n_10303), .Y (n_10305));
MX2X1 g31100(.A (n_6535), .B (n_6534), .S0 (n_10308), .Y (n_10309));
MX2X1 g31101(.A (n_6655), .B (n_6654), .S0 (n_10250), .Y (n_10307));
AOI22X1 g37723(.A0 (n_2558), .A1 (n_1242), .B0 (n_5516), .B1(n_1316), .Y (n_1243));
INVX1 g42298(.A (u9_mem_b2_b_116 ), .Y (n_2499));
NAND2X1 g39818(.A (u7_mem_b2_b_58 ), .B (n_12650), .Y (n_4116));
NAND2X1 g39819(.A (n_12389), .B (u4_mem_b0_b_102 ), .Y (n_11656));
NOR2X1 g30859(.A (n_10984), .B (n_11144), .Y (n_11146));
AOI21X1 g30858(.A0 (n_10615), .A1 (n_10196), .B0 (n_11144), .Y(n_11063));
NAND3X1 g30853(.A (n_9445), .B (n_1885), .C (n_8209), .Y (n_9545));
AOI21X1 g30852(.A0 (n_10621), .A1 (n_10202), .B0 (n_11069), .Y(n_11070));
AOI21X1 g30851(.A0 (n_10622), .A1 (n_10204), .B0 (n_5825), .Y(n_11072));
NAND3X1 g30850(.A (n_8844), .B (n_1886), .C (n_7530), .Y (n_9485));
AOI21X1 g30857(.A0 (n_10616), .A1 (n_10198), .B0 (n_11144), .Y(n_11064));
AOI21X1 g30856(.A0 (n_10618), .A1 (n_10199), .B0 (n_5825), .Y(n_11065));
AOI21X1 g30855(.A0 (n_10619), .A1 (n_10200), .B0 (n_11059), .Y(n_11066));
AOI21X1 g30854(.A0 (n_10620), .A1 (n_10201), .B0 (n_11144), .Y(n_11068));
INVX1 g42338(.A (u8_rp_b3_b ), .Y (n_494));
INVX1 g42335(.A (u11_mem_b3_b_57 ), .Y (n_6413));
INVX1 g42334(.A (u9_mem_b2_b_92 ), .Y (n_6902));
NOR2X1 g39915(.A (n_3089), .B (n_2744), .Y (n_2880));
NAND2X1 g39914(.A (u8_mem_b1_b_72 ), .B (n_12295), .Y (n_11456));
INVX2 g45498(.A (n_12076), .Y (n_12091));
AOI22X1 g37725(.A0 (n_6668), .A1 (n_2553), .B0 (n_6598), .B1(n_1316), .Y (n_2555));
NOR2X1 g39916(.A (n_3453), .B (n_2763), .Y (n_2879));
NAND2X1 g45948(.A (n_12334), .B (n_12336), .Y (n_12687));
NOR2X1 g39911(.A (n_3089), .B (n_2786), .Y (n_2883));
INVX1 g42567(.A (u11_mem_b3_b_67 ), .Y (n_6426));
NOR2X1 g39913(.A (n_3486), .B (n_2691), .Y (n_2882));
INVX1 g41575(.A (n_7443), .Y (n_675));
AOI22X1 g37726(.A0 (n_2558), .A1 (n_1685), .B0 (n_1684), .B1(n_1839), .Y (n_1686));
NOR2X1 g39912(.A (n_2681), .B (n_1488), .Y (n_1458));
NOR2X1 g39043(.A (n_2741), .B (n_1488), .Y (n_1423));
OR2X1 g41577(.A (n_1374), .B (n_5839), .Y (n_1375));
NAND2X1 g39734(.A (in_slt_415), .B (n_2368), .Y (n_4767));
MX2X1 g38620(.A (u4_mem_b0_b_91 ), .B (wb_din_661), .S0 (n_3765), .Y(n_3780));
NOR2X1 g40325(.A (n_1082), .B (n_2720), .Y (n_2666));
NAND2X1 g39737(.A (u5_mem_b2_b_34 ), .B (n_12823), .Y (n_12808));
INVX4 g41572(.A (n_743), .Y (n_5138));
CLKBUFX1 g45445(.A (n_12335), .Y (n_11827));
NAND2X1 g45943(.A (n_12684), .B (n_12685), .Y (n_12686));
NAND2X1 g39730(.A (n_3252), .B (u7_mem_b0_b_112 ), .Y (n_2993));
AOI21X1 g45942(.A0 (n_6317), .A1 (n_5751), .B0 (n_7214), .Y(n_12683));
INVX1 g39733(.A (n_4767), .Y (n_2989));
MX2X1 g38621(.A (u4_mem_b0_b_110 ), .B (wb_din_680), .S0 (n_3765), .Y(n_3779));
NAND2X1 g40795(.A (n_58), .B (u8_wp_b1_b ), .Y (n_937));
INVX2 g40794(.A (n_937), .Y (n_1129));
INVX1 g40791(.A (n_1129), .Y (n_2182));
AND2X1 g27(.A (n_9703), .B (n_9717), .Y (n_12589));
INVX1 g41853(.A (u7_rp_b3_b ), .Y (n_457));
CLKBUFX3 g45947(.A (n_12687), .Y (n_12688));
NOR2X1 g32907(.A (n_847), .B (o8_empty), .Y (n_9501));
NOR2X1 g32906(.A (n_12802), .B (o7_empty), .Y (n_9560));
NOR2X1 g32905(.A (n_12804), .B (o6_empty), .Y (n_9503));
NOR2X1 g32904(.A (n_854), .B (o4_empty), .Y (n_12846));
NOR2X1 g32903(.A (n_976), .B (o3_empty), .Y (n_12848));
NOR2X1 g32902(.A (n_9363), .B (n_10994), .Y (n_9517));
NAND2X1 g32901(.A (n_4633), .B (n_9513), .Y (n_9632));
INVX2 g32900(.A (n_9632), .Y (n_9675));
INVX1 g41857(.A (oc0_cfg_965), .Y (n_257));
INVX1 g41748(.A (n_829), .Y (n_1105));
NOR2X1 g32908(.A (n_977), .B (o9_empty), .Y (n_9499));
NAND2X1 g39106(.A (n_6044), .B (wb_addr_i_b4_b), .Y (n_1185));
NAND2X1 g39107(.A (n_2344), .B (in_slt_429), .Y (n_2357));
AOI21X1 g38072(.A0 (u8_mem_b3_b_146 ), .A1 (n_3879), .B0 (n_1498), .Y(n_3883));
INVX1 g41855(.A (oc4_cfg_1005), .Y (n_808));
INVX1 g41854(.A (n_808), .Y (n_4714));
NOR2X1 g39108(.A (n_4961), .B (n_2686), .Y (n_3446));
NOR2X1 g39109(.A (n_3453), .B (n_2804), .Y (n_3444));
NOR2X1 g40249(.A (n_995), .B (n_932), .Y (n_1224));
NOR2X1 g40248(.A (n_2477), .B (n_2864), .Y (n_2478));
MX2X1 g38623(.A (u4_mem_b0_b_112 ), .B (wb_din_682), .S0 (n_3765), .Y(n_3776));
NOR2X1 g40241(.A (n_867), .B (n_2712), .Y (n_2015));
NOR2X1 g40240(.A (n_935), .B (n_2829), .Y (n_2016));
NOR2X1 g40243(.A (n_2696), .B (n_3008), .Y (n_2697));
NOR2X1 g40242(.A (n_945), .B (n_2755), .Y (n_2014));
AOI21X1 g40245(.A0 (ic1_cfg_1034), .A1 (n_197), .B0(u14_u7_full_empty_r), .Y (n_974));
NOR2X1 g40244(.A (n_2041), .B (n_2765), .Y (n_2013));
NOR2X1 g40247(.A (n_2705), .B (n_2744), .Y (n_2694));
MX2X1 g36186(.A (n_6331), .B (n_6566), .S0 (n_6341), .Y (n_6332));
MX2X1 g38624(.A (u4_mem_b0_b_113 ), .B (wb_din_683), .S0 (n_3765), .Y(n_3773));
CLKBUFX3 g45962(.A (n_12738), .Y (n_12721));
INVX4 g45969(.A (n_12738), .Y (n_12735));
NOR2X1 g40309(.A (n_2477), .B (n_2763), .Y (n_1970));
NOR2X1 g40304(.A (n_2705), .B (n_2707), .Y (n_2673));
NOR2X1 g40305(.A (n_2093), .B (n_2782), .Y (n_1974));
NAND2X1 g40307(.A (n_5112), .B (n_4544), .Y (n_1972));
NOR2X1 g40300(.A (n_2736), .B (n_2801), .Y (n_2675));
NOR2X1 g40302(.A (n_935), .B (n_2732), .Y (n_1975));
NOR2X1 g40303(.A (n_1226), .B (n_2786), .Y (n_2674));
AOI21X1 g38059(.A0 (u3_mem_b3_b_151 ), .A1 (n_5138), .B0 (n_3392), .Y(n_5130));
AOI21X1 g38058(.A0 (u8_mem_b1_b_64 ), .A1 (n_4502), .B0 (n_1920), .Y(n_4503));
AOI21X1 g38053(.A0 (u3_mem_b3_b_138 ), .A1 (n_5138), .B0 (n_3151), .Y(n_5135));
AOI21X1 g38052(.A0 (u3_mem_b3_b_137 ), .A1 (n_5138), .B0 (n_2883), .Y(n_5136));
AOI21X1 g38051(.A0 (u3_mem_b3_b_136 ), .A1 (n_5133), .B0 (n_2851), .Y(n_5137));
AOI21X1 g38050(.A0 (u7_mem_b2_b_50 ), .A1 (n_4540), .B0 (n_2199), .Y(n_4506));
AOI21X1 g38057(.A0 (u3_mem_b3_b_144 ), .A1 (n_5138), .B0 (n_3400), .Y(n_5131));
AOI21X1 g38056(.A0 (u3_mem_b3_b_122 ), .A1 (n_5138), .B0 (n_3425), .Y(n_5132));
AOI21X1 g38055(.A0 (u3_mem_b3_b_140 ), .A1 (n_5133), .B0 (n_2905), .Y(n_5134));
AOI21X1 g38054(.A0 (u6_mem_b2_b_45 ), .A1 (n_4504), .B0 (n_2030), .Y(n_4505));
NOR2X1 g29976(.A (n_10809), .B (dma_ack_i_b1_b), .Y (n_11159));
NOR2X1 g29977(.A (n_10408), .B (dma_ack_i_b2_b), .Y (n_11124));
OR2X1 g29974(.A (u13_ints_r_b8_b ), .B (oc2_int_set), .Y (n_10830));
NOR2X1 g29975(.A (n_10409), .B (dma_ack_i_b0_b), .Y (n_11125));
OR2X1 g29973(.A (u13_ints_r_b5_b ), .B (oc1_int_set), .Y (n_10966));
OR2X1 g29971(.A (u13_ints_r_b17_b ), .B (oc5_int_set), .Y (n_10832));
NOR2X1 g29978(.A (n_10808), .B (dma_ack_i_b3_b), .Y (n_11158));
NOR2X1 g29979(.A (n_10407), .B (dma_ack_i_b4_b), .Y (n_11123));
AOI22X1 g37629(.A0 (n_6881), .A1 (n_1835), .B0 (n_6919), .B1(n_1760), .Y (n_1746));
AOI22X1 g37628(.A0 (n_2502), .A1 (n_6862), .B0 (n_6949), .B1(n_1859), .Y (n_1747));
OAI21X1 g37199(.A0 (u10_rp_b1_b ), .A1 (u10_wp_b2_b ), .B0 (n_480), .Y(n_1291));
XOR2X1 g37198(.A (n_798), .B (n_2594), .Y (n_2595));
XOR2X1 g37197(.A (n_1419), .B (n_4801), .Y (n_4802));
NAND2X1 g37194(.A (n_4617), .B (n_3416), .Y (n_6896));
NAND2X1 g37193(.A (n_4605), .B (n_3291), .Y (n_6925));
NAND2X1 g37192(.A (n_4098), .B (n_2238), .Y (n_6459));
NAND2X1 g37191(.A (n_2533), .B (n_2239), .Y (n_6003));
NAND2X1 g37190(.A (n_4555), .B (n_1796), .Y (n_6563));
OAI21X1 g33759(.A0 (n_4399), .A1 (n_9161), .B0 (n_7769), .Y (n_9121));
OAI21X1 g33758(.A0 (n_4323), .A1 (n_9161), .B0 (n_7770), .Y (n_9122));
OAI21X1 g33755(.A0 (n_4545), .A1 (n_9077), .B0 (n_7773), .Y (n_9127));
OAI21X1 g33754(.A0 (n_4543), .A1 (n_9110), .B0 (n_7774), .Y (n_9128));
OAI21X1 g33757(.A0 (n_4358), .A1 (n_9139), .B0 (n_7771), .Y (n_9124));
OAI21X1 g33756(.A0 (n_4547), .A1 (n_9170), .B0 (n_7772), .Y (n_9125));
OAI21X1 g33751(.A0 (n_4334), .A1 (n_9161), .B0 (n_7777), .Y (n_9131));
OAI21X1 g33750(.A0 (n_4535), .A1 (n_9182), .B0 (n_7778), .Y (n_9132));
OAI21X1 g33753(.A0 (n_4332), .A1 (n_9139), .B0 (n_7775), .Y (n_9129));
OAI21X1 g33752(.A0 (n_4539), .A1 (n_9139), .B0 (n_7776), .Y (n_9130));
AOI21X1 g37997(.A0 (u6_mem_b2_b_54 ), .A1 (n_4504), .B0 (n_2162), .Y(n_4543));
AOI21X1 g37996(.A0 (u3_mem_b1_b_89 ), .A1 (n_5157), .B0 (n_2655), .Y(n_5156));
NOR2X1 g35856(.A (n_2625), .B (n_4851), .Y (n_4852));
AOI21X1 g37994(.A0 (u7_mem_b2_b_31 ), .A1 (n_4540), .B0 (n_2021), .Y(n_4546));
AOI21X1 g37993(.A0 (u3_mem_b1_b_61 ), .A1 (n_5157), .B0 (n_2662), .Y(n_5158));
AOI21X1 g37992(.A0 (u7_mem_b3_b_141 ), .A1 (n_5145), .B0 (n_3407), .Y(n_5159));
AOI21X1 g37991(.A0 (u6_mem_b2_b_56 ), .A1 (n_4544), .B0 (n_2223), .Y(n_4547));
AOI21X1 g37990(.A0 (u3_mem_b1_b_87 ), .A1 (n_5157), .B0 (n_2769), .Y(n_5160));
INVX2 g40872(.A (n_1430), .Y (n_2705));
BUFX3 g40871(.A (n_1226), .Y (n_5069));
INVX2 g40876(.A (n_1226), .Y (n_1430));
INVX1 g40877(.A (n_1430), .Y (n_2721));
AOI21X1 g37999(.A0 (u5_mem_b2_b_41 ), .A1 (n_4378), .B0 (n_1838), .Y(n_4542));
AOI21X1 g37998(.A0 (u3_mem_b1_b_90 ), .A1 (n_5157), .B0 (n_2728), .Y(n_5155));
NAND2X1 g37448(.A (u13_ints_r_b10_b ), .B (n_3979), .Y (n_3981));
INVX2 g33285(.A (n_12689), .Y (n_10605));
AOI21X1 g33284(.A0 (n_7157), .A1 (n_1230), .B0 (n_7434), .Y (n_7387));
AOI21X1 g33283(.A0 (n_7031), .A1 (n_1105), .B0 (n_7378), .Y (n_7294));
AOI21X1 g33282(.A0 (n_7032), .A1 (n_1136), .B0 (n_7379), .Y (n_7295));
NAND3X1 g33281(.A (n_9833), .B (n_657), .C (n_7870), .Y (n_8178));
NAND2X1 g33280(.A (n_9710), .B (u15_crac_rd), .Y (n_9882));
BUFX3 g37441(.A (n_7297), .Y (n_7468));
AOI21X1 g38216(.A0 (u7_mem_b1_b_67 ), .A1 (n_5118), .B0 (n_2807), .Y(n_5079));
NAND2X1 g37445(.A (n_2575), .B (n_838), .Y (n_2588));
INVX2 g37444(.A (n_2588), .Y (n_7297));
NAND2X1 g37447(.A (u13_ints_r_b0_b ), .B (n_3979), .Y (n_3982));
NAND3X1 g37446(.A (n_593), .B (n_7443), .C (n_2574), .Y (n_2587));
AOI21X1 g45863(.A0 (n_12588), .A1 (n_12589), .B0 (n_12590), .Y(n_12591));
INVX1 g42516(.A (u11_mem_b0_b_159 ), .Y (n_6372));
OAI21X1 g35858(.A0 (n_5701), .A1 (n_11934), .B0 (n_6238), .Y(n_7105));
NAND2X1 g31667(.A (n_1748), .B (n_10073), .Y (n_9991));
NAND2X1 g31666(.A (n_337), .B (n_10081), .Y (n_9992));
NAND2X1 g31665(.A (n_312), .B (n_10391), .Y (n_10392));
NAND2X1 g31664(.A (n_334), .B (n_10391), .Y (n_10393));
NAND2X1 g31663(.A (n_314), .B (n_10081), .Y (n_9993));
OR2X1 g31662(.A (n_9497), .B (n_9486), .Y (n_9612));
OR2X1 g31661(.A (n_9559), .B (n_9548), .Y (n_9660));
OR2X1 g31660(.A (n_9498), .B (n_9488), .Y (n_9615));
NOR2X1 g45682(.A (n_11673), .B (dma_ack_i_b7_b), .Y (n_12379));
INVX1 g42651(.A (oc2_int_set_712), .Y (n_450));
INVX1 g42652(.A (u11_mem_b1_b_146 ), .Y (n_1595));
INVX1 g42653(.A (u9_mem_b2_b_89 ), .Y (n_6933));
NOR2X1 g31669(.A (n_11892), .B (n_11586), .Y (n_9990));
OR2X1 g31668(.A (n_9558), .B (n_9546), .Y (n_9657));
NAND2X1 g39483(.A (n_1225), .B (n_1300), .Y (n_1271));
INVX1 g39480(.A (n_1271), .Y (n_4729));
NAND2X1 g39487(.A (n_12204), .B (u6_mem_b0_b_94 ), .Y (n_11709));
NAND2X1 g39486(.A (u4_mem_b1_b_83 ), .B (n_12265), .Y (n_4183));
NAND2X1 g39485(.A (n_12721), .B (u3_mem_b0_b_93 ), .Y (n_3150));
NOR2X1 g39484(.A (n_5138), .B (n_2735), .Y (n_3151));
INVX8 g35108(.A (o6_we), .Y (n_7870));
NAND2X1 g39488(.A (u8_mem_b2_b_33 ), .B (n_2362), .Y (n_2295));
MX2X1 g36716(.A (u10_mem_b2_b_106 ), .B (n_5422), .S0 (n_5424), .Y(n_5425));
AOI21X1 g36717(.A0 (n_5580), .A1 (n_6649), .B0 (n_4804), .Y (n_5581));
AOI21X1 g36714(.A0 (n_5582), .A1 (n_6649), .B0 (n_4803), .Y (n_5583));
MX2X1 g36715(.A (u10_mem_b2_b_105 ), .B (n_5418), .S0 (n_5424), .Y(n_5426));
OAI21X1 g36712(.A0 (n_4571), .A1 (n_5169), .B0 (n_6152), .Y (n_5742));
MX2X1 g36713(.A (u11_mem_b0_b_167 ), .B (n_5413), .S0 (n_6359), .Y(n_5428));
OAI21X1 g36710(.A0 (n_4551), .A1 (n_5161), .B0 (n_6152), .Y (n_5743));
NAND2X1 g36711(.A (n_5559), .B (n_6091), .Y (n_6092));
CLKBUFX3 g45541(.A (n_12148), .Y (n_12149));
MX2X1 g36718(.A (u9_mem_b0_b_167 ), .B (n_5736), .S0 (n_6856), .Y(n_5740));
MX2X1 g36719(.A (u9_mem_b0_b_168 ), .B (n_5733), .S0 (n_6856), .Y(n_5738));
INVX1 g42436(.A (u11_mem_b0_b_163 ), .Y (n_6363));
INVX1 g42437(.A (u10_mem_b0_b ), .Y (n_5959));
INVX1 g42430(.A (u11_mem_b2_b_115 ), .Y (n_188));
NAND2X1 g32743(.A (n_341), .B (n_10605), .Y (n_12017));
INVX1 g42432(.A (u10_mem_b2_b_110 ), .Y (n_366));
NOR2X1 g45542(.A (u14_u1_en_out_l2), .B (n_8670), .Y (n_12148));
INVX1 g42438(.A (u11_mem_b2_b_91 ), .Y (n_6439));
NAND2X1 g31591(.A (n_1679), .B (n_10054), .Y (n_10062));
NAND2X1 g31590(.A (n_356), .B (n_10054), .Y (n_10063));
NAND2X1 g31593(.A (n_340), .B (n_10054), .Y (n_10059));
NAND2X1 g31592(.A (n_1737), .B (n_10054), .Y (n_10060));
NAND2X1 g31595(.A (n_45), .B (n_10054), .Y (n_10057));
NAND2X1 g31594(.A (n_42), .B (n_10010), .Y (n_10058));
NAND2X1 g31597(.A (n_1727), .B (n_10054), .Y (n_10055));
NAND2X1 g31596(.A (n_1703), .B (n_10054), .Y (n_10056));
NAND2X1 g31599(.A (n_206), .B (n_10054), .Y (n_10052));
NAND2X1 g31598(.A (n_1723), .B (n_10054), .Y (n_10053));
INVX2 g40494(.A (wb_din_685), .Y (n_2831));
OAI21X1 g45549(.A0 (n_5542), .A1 (n_7080), .B0 (n_6200), .Y(n_12157));
NOR2X1 g39664(.A (n_3117), .B (n_2744), .Y (n_3027));
NAND2X1 g39663(.A (n_2302), .B (in_slt_422), .Y (n_2268));
NAND2X1 g39660(.A (n_2325), .B (in_slt_450), .Y (n_2269));
NAND2X1 g36909(.A (n_2540), .B (n_2537), .Y (n_4815));
NAND4X1 g36908(.A (n_12841), .B (n_12842), .C (n_12041), .D (n_1333),.Y (n_5561));
NAND4X1 g36902(.A (n_12855), .B (n_12856), .C (n_12798), .D (n_1534),.Y (n_5879));
INVX2 g36906(.A (n_5561), .Y (n_5562));
NAND4X1 g36905(.A (n_12805), .B (n_12806), .C (n_3229), .D (n_1541),.Y (n_5713));
NAND2X1 g38992(.A (u7_mem_b3_b_126 ), .B (n_1538), .Y (n_1506));
NAND2X1 g36421(.A (n_5898), .B (n_6259), .Y (n_5899));
NAND2X1 g37545(.A (n_554), .B (in_slt_742), .Y (n_1007));
MX2X1 g33993(.A (u4_mem_b0_b_110 ), .B (n_3779), .S0 (n_7499), .Y(n_8827));
MX2X1 g33992(.A (u4_mem_b0_b_91 ), .B (n_3780), .S0 (n_7499), .Y(n_8829));
MX2X1 g33991(.A (u4_mem_b0_b_109 ), .B (n_3783), .S0 (n_7499), .Y(n_9439));
MX2X1 g33990(.A (u4_mem_b0_b_108 ), .B (n_3784), .S0 (n_7499), .Y(n_8830));
MX2X1 g33997(.A (u4_mem_b0_b_114 ), .B (n_3770), .S0 (n_7499), .Y(n_9435));
MX2X1 g33996(.A (u4_mem_b0_b_113 ), .B (n_3773), .S0 (n_7499), .Y(n_8824));
MX2X1 g33995(.A (u4_mem_b0_b_112 ), .B (n_3776), .S0 (n_7499), .Y(n_9437));
MX2X1 g33994(.A (u4_mem_b0_b_111 ), .B (n_3777), .S0 (n_7499), .Y(n_8825));
MX2X1 g38742(.A (u3_mem_b0_b_91 ), .B (wb_din_661), .S0 (n_3807), .Y(n_3598));
MX2X1 g33999(.A (u4_mem_b0_b_116 ), .B (n_3766), .S0 (n_7499), .Y(n_8822));
MX2X1 g33998(.A (u4_mem_b0_b_115 ), .B (n_3768), .S0 (n_7499), .Y(n_8823));
OAI21X1 g33903(.A0 (n_4877), .A1 (n_8948), .B0 (n_7620), .Y (n_8944));
AOI21X1 g38572(.A0 (u3_mem_b1_b_81 ), .A1 (n_5148), .B0 (n_2658), .Y(n_4860));
MX2X1 g38740(.A (u8_mem_b0_b_104 ), .B (wb_din_674), .S0 (n_3826), .Y(n_3600));
NAND2X1 g34419(.A (u4_mem_b2_b_57 ), .B (n_7984), .Y (n_7997));
NAND2X1 g34418(.A (u4_mem_b2_b_56 ), .B (n_7984), .Y (n_7998));
NAND2X1 g34417(.A (u4_mem_b2_b_55 ), .B (n_7984), .Y (n_7999));
NAND2X1 g34416(.A (u4_mem_b2_b_54 ), .B (n_7984), .Y (n_8000));
NAND2X1 g34415(.A (u4_mem_b2_b_53 ), .B (n_7984), .Y (n_8001));
NAND2X1 g34414(.A (n_7444), .B (n_996), .Y (n_7518));
MX2X1 g38747(.A (u8_mem_b0_b_115 ), .B (wb_din_685), .S0 (n_3826), .Y(n_3590));
NAND2X1 g38993(.A (u8_mem_b3_b_145 ), .B (n_2468), .Y (n_2375));
AOI21X1 g38443(.A0 (u6_mem_b3_b_136 ), .A1 (n_5059), .B0 (n_3410), .Y(n_4923));
MX2X1 g38746(.A (u3_mem_b0_b_113 ), .B (wb_din_683), .S0 (n_3807), .Y(n_3592));
AOI21X1 g38444(.A0 (u4_mem_b2_b_48 ), .A1 (n_935), .B0 (n_1975), .Y(n_4327));
MX2X1 g38745(.A (u3_mem_b0_b_111 ), .B (wb_din_681), .S0 (n_3807), .Y(n_3593));
XOR2X1 g40403(.A (n_7048), .B (n_888), .Y (n_1806));
INVX8 g41754(.A (n_1103), .Y (n_3765));
NAND2X1 g32718(.A (n_157), .B (n_10605), .Y (n_11750));
NAND2X1 g32719(.A (n_195), .B (n_10605), .Y (n_11724));
NAND2X1 g32712(.A (n_362), .B (n_10617), .Y (n_10609));
NAND2X1 g32713(.A (n_376), .B (n_10617), .Y (n_12794));
NAND2X1 g32710(.A (n_280), .B (n_10617), .Y (n_12196));
NAND2X1 g32711(.A (n_352), .B (n_10617), .Y (n_12065));
NAND2X1 g32716(.A (n_389), .B (n_10605), .Y (n_11744));
NAND2X1 g32717(.A (n_398), .B (n_10605), .Y (n_11746));
NAND2X1 g32714(.A (n_384), .B (n_10617), .Y (n_10607));
NAND2X1 g32715(.A (n_12688), .B (n_862), .Y (n_11099));
AOI21X1 g38422(.A0 (u6_mem_b2_b_38 ), .A1 (n_4504), .B0 (n_2080), .Y(n_4338));
AOI21X1 g38423(.A0 (u7_mem_b1_b_78 ), .A1 (n_5069), .B0 (n_2693), .Y(n_4932));
AOI21X1 g38420(.A0 (u6_mem_b1_b_65 ), .A1 (n_5019), .B0 (n_2727), .Y(n_4934));
AOI21X1 g38421(.A0 (u6_mem_b1_b_71 ), .A1 (n_5112), .B0 (n_2838), .Y(n_4933));
AOI21X1 g38426(.A0 (u6_mem_b2_b_44 ), .A1 (n_4504), .B0 (n_2190), .Y(n_4336));
AOI21X1 g38427(.A0 (u7_mem_b3_b_126 ), .A1 (n_4961), .B0 (n_3032), .Y(n_4931));
AOI21X1 g38424(.A0 (u8_mem_b3_b_150 ), .A1 (n_3879), .B0 (n_1273), .Y(n_3854));
AOI21X1 g38425(.A0 (u6_mem_b2_b_42 ), .A1 (n_4504), .B0 (n_1968), .Y(n_4337));
NOR2X1 g39418(.A (u10_mem_b1_b_137 ), .B (n_2364), .Y (n_2307));
AOI21X1 g38428(.A0 (u6_mem_b2_b_29 ), .A1 (n_4504), .B0 (n_1996), .Y(n_4335));
AOI21X1 g38429(.A0 (u6_mem_b1_b_69 ), .A1 (n_5019), .B0 (n_2676), .Y(n_4930));
OAI21X1 g30904(.A0 (n_7294), .A1 (n_7524), .B0 (n_8909), .Y (n_9473));
INVX1 g33300(.A (n_12149), .Y (n_9947));
INVX2 g41021(.A (n_7080), .Y (n_6773));
OAI21X1 g33805(.A0 (n_4867), .A1 (n_8393), .B0 (n_7589), .Y (n_9067));
NAND2X1 g34272(.A (u3_mem_b2_b_47 ), .B (n_8141), .Y (n_8127));
OAI21X1 g33807(.A0 (n_4905), .A1 (n_9034), .B0 (n_7721), .Y (n_9065));
OAI21X1 g33806(.A0 (n_4902), .A1 (n_9034), .B0 (n_7722), .Y (n_9066));
MX2X1 g37298(.A (u11_mem_b2_b_113 ), .B (n_5309), .S0 (n_5312), .Y(n_5310));
MX2X1 g37299(.A (u11_mem_b2_b_114 ), .B (n_5307), .S0 (n_5312), .Y(n_5308));
MX2X1 g37294(.A (u11_mem_b2_b_108 ), .B (n_5317), .S0 (n_5409), .Y(n_5318));
OAI21X1 g33801(.A0 (n_4343), .A1 (n_8440), .B0 (n_8122), .Y (n_9071));
MX2X1 g37296(.A (u11_mem_b2_b_110 ), .B (n_5313), .S0 (n_5312), .Y(n_5314));
MX2X1 g37297(.A (u11_mem_b2_b_112 ), .B (n_5280), .S0 (n_5312), .Y(n_5311));
MX2X1 g37290(.A (u11_mem_b1_b_139 ), .B (n_5317), .S0 (n_6502), .Y(n_5323));
MX2X1 g37291(.A (u11_mem_b2_b_111 ), .B (n_5321), .S0 (n_5409), .Y(n_5322));
MX2X1 g37292(.A (u11_mem_b1_b_146 ), .B (n_5304), .S0 (n_5405), .Y(n_5320));
OAI21X1 g33556(.A0 (n_4423), .A1 (n_8333), .B0 (n_8001), .Y (n_8282));
NAND2X1 g36479(.A (n_5869), .B (n_1229), .Y (n_5870));
NAND2X1 g36478(.A (n_5874), .B (n_5876), .Y (n_5871));
OAI21X1 g33555(.A0 (n_4425), .A1 (n_8333), .B0 (n_8002), .Y (n_8283));
OAI21X1 g33802(.A0 (n_3852), .A1 (n_8438), .B0 (n_8134), .Y (n_9070));
NAND2X1 g36477(.A (n_12681), .B (n_6141), .Y (n_5873));
NOR2X1 g36476(.A (n_2609), .B (n_1776), .Y (n_5440));
INVX2 g36475(.A (n_5440), .Y (n_11119));
OAI21X1 g33908(.A0 (n_4388), .A1 (n_8449), .B0 (n_7948), .Y (n_8938));
NAND2X1 g34279(.A (u3_mem_b2_b_54 ), .B (n_8101), .Y (n_8121));
BUFX3 g40710(.A (n_941), .Y (n_4544));
MX2X1 g38725(.A (u7_mem_b0_b_93 ), .B (wb_din_663), .S0 (n_3622), .Y(n_3616));
OAI21X1 g33904(.A0 (n_4484), .A1 (n_8856), .B0 (n_7617), .Y (n_8943));
NAND2X1 g34625(.A (u6_mem_b1_b_62 ), .B (n_7758), .Y (n_7800));
NAND2X1 g36338(.A (n_5865), .B (n_3559), .Y (n_5929));
NAND2X1 g34626(.A (u6_mem_b1_b_63 ), .B (n_7758), .Y (n_7799));
NAND2X1 g36339(.A (n_6248), .B (n_6824), .Y (n_6313));
NAND2X1 g34627(.A (u6_mem_b1_b_64 ), .B (n_7758), .Y (n_7798));
NAND2X1 g34620(.A (u8_mem_b2_b_39 ), .B (n_7976), .Y (n_7805));
MX2X1 g38724(.A (u6_mem_b0_b_117 ), .B (wb_din_687), .S0 (n_3632), .Y(n_3617));
NAND2X1 g34621(.A (u6_mem_b1_b_88 ), .B (n_7758), .Y (n_7804));
NAND2X1 g34622(.A (u6_mem_b1_b_61 ), .B (n_7758), .Y (n_7803));
NAND2X1 g34623(.A (u6_mem_b1_b_89 ), .B (n_7758), .Y (n_7802));
NAND2X1 g37870(.A (n_4150), .B (n_3472), .Y (n_12058));
AOI22X1 g37871(.A0 (n_5969), .A1 (n_1575), .B0 (n_6035), .B1(n_1831), .Y (n_1566));
NAND2X1 g37872(.A (n_2400), .B (n_3084), .Y (n_4574));
NAND2X1 g37873(.A (n_4244), .B (n_3057), .Y (n_5200));
AOI22X1 g37874(.A0 (u10_din_tmp_53), .A1 (n_3339), .B0 (n_3911), .B1(in_slt_432), .Y (n_3910));
NAND2X1 g37875(.A (n_2462), .B (n_3054), .Y (n_4573));
NAND2X1 g37876(.A (n_4159), .B (n_3519), .Y (n_5199));
NAND2X1 g37877(.A (n_2418), .B (n_3051), .Y (n_4572));
NAND2X1 g37878(.A (n_4212), .B (n_2995), .Y (n_5198));
AOI22X1 g37879(.A0 (u10_din_tmp_54), .A1 (n_3339), .B0 (n_3911), .B1(in_slt_433), .Y (n_3909));
MX2X1 g33141(.A (wb_din_673), .B (n_8565), .S0 (n_8538), .Y (n_8566));
MX2X1 g33142(.A (wb_din_674), .B (oc1_cfg_979), .S0 (n_8538), .Y(n_8564));
MX2X1 g33143(.A (wb_din_675), .B (oc1_cfg_980), .S0 (n_8538), .Y(n_8563));
MX2X1 g33144(.A (wb_din_676), .B (n_9833), .S0 (n_8538), .Y (n_8562));
MX2X1 g33146(.A (wb_din_678), .B (oc2_cfg_985), .S0 (n_8538), .Y(n_8558));
MX2X1 g33147(.A (wb_din_679), .B (oc2_cfg_986), .S0 (n_8538), .Y(n_8556));
MX2X1 g33148(.A (wb_din_661), .B (oc0_cfg_964), .S0 (n_8538), .Y(n_8555));
MX2X1 g33149(.A (wb_din_680), .B (oc2_cfg_987), .S0 (n_8538), .Y(n_8554));
INVX8 g41513(.A (n_1076), .Y (n_3807));
INVX2 g41511(.A (n_858), .Y (n_1076));
MX2X1 g36114(.A (n_6445), .B (n_6444), .S0 (n_5312), .Y (n_6446));
MX2X1 g38726(.A (u6_mem_b0_b_115 ), .B (wb_din_685), .S0 (n_3632), .Y(n_3615));
NAND2X1 g36443(.A (n_6248), .B (n_12531), .Y (n_6249));
NAND2X1 g36440(.A (n_6250), .B (n_1038), .Y (n_6251));
MX2X1 g31128(.A (n_6889), .B (n_6888), .S0 (n_10277), .Y (n_10272));
MX2X1 g31129(.A (n_6932), .B (n_6931), .S0 (n_10235), .Y (n_10270));
MX2X1 g36117(.A (n_6437), .B (n_6544), .S0 (n_5312), .Y (n_6438));
MX2X1 g31120(.A (n_6639), .B (n_6638), .S0 (n_10267), .Y (n_10283));
MX2X1 g31121(.A (n_6636), .B (n_6635), .S0 (n_10267), .Y (n_10281));
MX2X1 g31122(.A (n_6874), .B (n_6873), .S0 (n_10267), .Y (n_10280));
MX2X1 g31123(.A (n_6936), .B (n_6935), .S0 (n_10277), .Y (n_10279));
MX2X1 g31124(.A (n_6882), .B (n_6881), .S0 (n_10277), .Y (n_10278));
MX2X1 g31125(.A (n_6634), .B (n_6633), .S0 (n_10137), .Y (n_10276));
MX2X1 g31126(.A (n_6934), .B (n_6933), .S0 (n_10277), .Y (n_10275));
MX2X1 g31127(.A (n_6631), .B (n_6630), .S0 (n_10137), .Y (n_10274));
NAND2X1 g39872(.A (u4_mem_b1_b_86 ), .B (n_12270), .Y (n_4112));
NAND2X1 g39873(.A (n_12679), .B (u5_mem_b0_b_111 ), .Y (n_3840));
NAND2X1 g39870(.A (n_2344), .B (in_slt4), .Y (n_2236));
NAND2X1 g39871(.A (n_1205), .B (u5_rp_b3_b ), .Y (n_4644));
NAND2X1 g39876(.A (n_2491), .B (u7_mem_b0_b_119 ), .Y (n_2479));
NAND2X1 g39877(.A (u3_mem_b2_b_52 ), .B (n_3330), .Y (n_2636));
NOR2X1 g39874(.A (n_3453), .B (n_2702), .Y (n_2909));
NAND2X1 g39875(.A (u6_mem_b2_b_50 ), .B (n_3423), .Y (n_2908));
NAND2X1 g39878(.A (u6_mem_b2_b_34 ), .B (n_2285), .Y (n_2482));
NAND2X1 g36445(.A (n_3940), .B (n_5466), .Y (n_7010));
NAND2X1 g31645(.A (n_5504), .B (n_10010), .Y (n_9999));
NOR2X1 g45881(.A (n_11533), .B (n_8667), .Y (n_12607));
NAND2X1 g31644(.A (n_5506), .B (n_10010), .Y (n_10000));
NAND2X1 g31647(.A (n_10992), .B (u4_rp_b0_b ), .Y (n_9843));
AOI22X1 g37707(.A0 (n_2558), .A1 (n_5949), .B0 (n_6028), .B1(n_2544), .Y (n_1687));
INVX1 g42358(.A (u9_mem_b3_b_75 ), .Y (n_6087));
MX2X1 g38720(.A (u7_mem_b0_b_97 ), .B (wb_din_667), .S0 (n_3622), .Y(n_3623));
NAND3X1 g31646(.A (n_9641), .B (n_11600), .C (n_9564), .Y (n_9844));
INVX1 g42353(.A (in_slt_738), .Y (n_197));
INVX1 g42352(.A (u6_rp_b3_b ), .Y (n_496));
INVX1 g42355(.A (u11_mem_b0_b_153 ), .Y (n_6353));
INVX1 g42354(.A (u10_mem_b3_b_64 ), .Y (n_6002));
INVX1 g42357(.A (oc5_cfg_1016), .Y (n_127));
NAND2X1 g31640(.A (n_5359), .B (n_10065), .Y (n_10004));
NAND2X1 g38984(.A (u5_mem_b3_b_142 ), .B (n_3543), .Y (n_3527));
NOR2X1 g35817(.A (n_453), .B (n_6752), .Y (n_6753));
NAND2X1 g31643(.A (n_5510), .B (n_10010), .Y (n_10001));
MX2X1 g38723(.A (u7_mem_b0_b_94 ), .B (wb_din_664), .S0 (n_3622), .Y(n_3619));
AOI22X1 g37823(.A0 (n_1756), .A1 (n_1610), .B0 (n_1609), .B1(n_1643), .Y (n_1611));
NAND2X1 g38987(.A (u3_mem_b3_b_138 ), .B (n_1517), .Y (n_1508));
MX2X1 g38722(.A (u7_mem_b0_b_95 ), .B (wb_din_665), .S0 (n_3622), .Y(n_3620));
MX2X1 g38718(.A (u7_mem_b0_b_98 ), .B (wb_din_668), .S0 (n_3622), .Y(n_3625));
MX2X1 g38719(.A (u5_mem_b0_b_103 ), .B (wb_din_673), .S0 (n_3720), .Y(n_3624));
AOI21X1 g31657(.A0 (n_7165), .A1 (n_1071), .B0 (n_9560), .Y (n_9561));
AND2X1 g38986(.A (n_996), .B (n_1300), .Y (n_1132));
NOR2X1 g39296(.A (n_3486), .B (n_2755), .Y (n_3844));
NOR2X1 g39297(.A (n_3486), .B (n_2741), .Y (n_3305));
NOR2X1 g39294(.A (n_3486), .B (n_2681), .Y (n_3307));
NOR2X1 g39292(.A (n_5102), .B (n_2829), .Y (n_3309));
NOR2X1 g39293(.A (u10_mem_b1_b_141 ), .B (n_2364), .Y (n_2327));
NAND2X1 g39290(.A (n_12204), .B (u6_mem_b0_b_101 ), .Y (n_11707));
NOR2X1 g39291(.A (n_3453), .B (n_2691), .Y (n_3311));
NOR2X1 g39298(.A (n_3486), .B (n_2735), .Y (n_3302));
AOI21X1 g45544(.A0 (n_12152), .A1 (n_12153), .B0 (n_12640), .Y(n_12156));
MX2X1 g38608(.A (u4_mem_b0_b_101 ), .B (wb_din_671), .S0 (n_3765), .Y(n_3801));
NOR2X1 g35812(.A (n_597), .B (n_5440), .Y (n_6741));
MX2X1 g38710(.A (u7_mem_b0_b_118 ), .B (wb_din_688), .S0 (n_3622), .Y(n_3636));
INVX4 g32960(.A (n_10376), .Y (n_9903));
NAND2X1 g32963(.A (n_3944), .B (n_9571), .Y (n_9674));
INVX2 g32962(.A (n_9674), .Y (n_9720));
NOR2X1 g32965(.A (o4_empty), .B (n_458), .Y (n_9559));
NOR2X1 g32964(.A (o3_empty), .B (n_459), .Y (n_9498));
NOR2X1 g32967(.A (o7_empty), .B (n_422), .Y (n_9558));
NOR2X1 g32966(.A (o6_empty), .B (n_447), .Y (n_9497));
AND2X1 g32969(.A (n_9705), .B (n_9719), .Y (n_11131));
INVX1 g32968(.A (n_11131), .Y (n_9902));
AND2X1 g36642(.A (n_3973), .B (n_4733), .Y (n_5585));
INVX1 g43009(.A (n_1036), .Y (n_715));
NAND2X1 g39120(.A (u6_mem_b1_b_86 ), .B (n_12169), .Y (n_4229));
NAND2X1 g39121(.A (u4_mem_b2_b_36 ), .B (n_12079), .Y (n_2355));
NOR2X1 g40261(.A (n_2741), .B (n_1985), .Y (n_1884));
NOR2X1 g40260(.A (n_2782), .B (n_1985), .Y (n_2002));
NOR2X1 g39124(.A (n_3486), .B (n_2786), .Y (n_3434));
INVX1 g37076(.A (n_12116), .Y (n_5680));
OR2X1 g39126(.A (n_3431), .B (n_1200), .Y (n_3432));
NOR2X1 g40264(.A (n_2470), .B (n_2765), .Y (n_2481));
NOR2X1 g40269(.A (n_2470), .B (n_2804), .Y (n_2483));
NOR2X1 g40268(.A (n_935), .B (n_2790), .Y (n_1998));
AOI22X1 g37827(.A0 (n_298), .A1 (n_1575), .B0 (n_5500), .B1 (n_1831),.Y (n_1603));
NAND2X1 g36643(.A (n_5279), .B (n_3981), .Y (n_5786));
NOR2X1 g40062(.A (n_2794), .B (n_1985), .Y (n_2165));
AOI22X1 g37826(.A0 (n_1756), .A1 (n_1605), .B0 (n_1604), .B1(n_1643), .Y (n_1606));
MX2X1 g38607(.A (u4_mem_b0_b_100 ), .B (wb_din_670), .S0 (n_3765), .Y(n_3802));
AOI21X1 g40067(.A0 (oc3_cfg_994), .A1 (in_slt_749), .B0(u14_u3_full_empty_r), .Y (n_553));
NAND2X1 g34489(.A (u5_mem_b1_b ), .B (n_7870), .Y (n_7943));
NAND2X1 g45985(.A (n_656), .B (n_601), .Y (n_12751));
INVX2 g45984(.A (n_12751), .Y (n_12752));
NAND2X1 g45981(.A (u3_mem_b3_b_135 ), .B (n_2463), .Y (n_12750));
NAND2X1 g45980(.A (n_3207), .B (u3_mem_b2_b_42 ), .Y (n_12749));
CLKBUFX1 g45983(.A (n_12752), .Y (n_12753));
NAND2X2 g45982(.A (n_12753), .B (u3_mem_b1_b_73 ), .Y (n_12754));
AOI22X1 g37825(.A0 (n_2558), .A1 (n_5962), .B0 (n_6037), .B1 (n_940),.Y (n_2525));
MX2X1 g34066(.A (u6_mem_b0_b_117 ), .B (n_3617), .S0 (n_7505), .Y(n_8764));
MX2X1 g34067(.A (u6_mem_b0_b_118 ), .B (n_3621), .S0 (n_7505), .Y(n_8763));
MX2X1 g34064(.A (u6_mem_b0_b_115 ), .B (n_3615), .S0 (n_7505), .Y(n_8766));
MX2X1 g34065(.A (u6_mem_b0_b_116 ), .B (n_3670), .S0 (n_7505), .Y(n_8765));
MX2X1 g34062(.A (u6_mem_b0_b_113 ), .B (n_3671), .S0 (n_7505), .Y(n_8767));
MX2X1 g34063(.A (u6_mem_b0_b_114 ), .B (n_3614), .S0 (n_7505), .Y(n_9407));
MX2X1 g34060(.A (u6_mem_b0_b_111 ), .B (n_3608), .S0 (n_7505), .Y(n_8768));
MX2X1 g34061(.A (u6_mem_b0_b_112 ), .B (n_3611), .S0 (n_7505), .Y(n_9409));
NAND2X1 g38923(.A (u4_mem_b3_b_141 ), .B (n_3556), .Y (n_3531));
MX2X1 g34068(.A (u6_mem_b0_b_119 ), .B (n_3633), .S0 (n_7505), .Y(n_8761));
MX2X1 g34069(.A (u6_mem_b0_b_92 ), .B (n_3668), .S0 (n_7505), .Y(n_8760));
OAI21X1 g33817(.A0 (n_4932), .A1 (n_9055), .B0 (n_7708), .Y (n_9050));
AOI22X1 g37824(.A0 (n_270), .A1 (n_1575), .B0 (n_5492), .B1 (n_1831),.Y (n_1607));
MX2X1 g38605(.A (u3_mem_b0_b_105 ), .B (wb_din_675), .S0 (n_3807), .Y(n_3804));
NAND2X1 g38922(.A (u4_mem_b3_b_131 ), .B (n_3546), .Y (n_3532));
NAND2X1 g39180(.A (n_12389), .B (u4_mem_b0_b_108 ), .Y (n_2972));
AOI21X1 g38398(.A0 (u3_mem_b2_b_55 ), .A1 (n_4519), .B0 (n_1955), .Y(n_4341));
AND2X1 g34487(.A (n_7286), .B (n_7443), .Y (n_7514));
NAND2X1 g38921(.A (u5_mem_b3_b_146 ), .B (n_3543), .Y (n_2401));
AND2X1 g29952(.A (n_10967), .B (n_11119), .Y (n_11121));
AND2X1 g29953(.A (n_10833), .B (n_11119), .Y (n_11015));
AND2X1 g29954(.A (n_10832), .B (n_11119), .Y (n_11014));
AND2X1 g29955(.A (n_10831), .B (n_11119), .Y (n_11012));
AND2X1 g29956(.A (n_10966), .B (n_11119), .Y (n_11120));
AND2X1 g29957(.A (n_10830), .B (n_11119), .Y (n_11011));
NAND2X1 g37607(.A (n_3521), .B (n_3436), .Y (n_4631));
NAND2X1 g37606(.A (n_3554), .B (n_3497), .Y (n_4632));
AOI22X1 g37605(.A0 (n_785), .A1 (n_3543), .B0 (n_3559), .B1(u5_rp_b3_b ), .Y (n_3939));
AOI22X1 g37604(.A0 (n_650), .A1 (n_1546), .B0 (n_12634), .B1(u7_rp_b3_b ), .Y (n_1772));
AOI22X1 g37603(.A0 (n_664), .A1 (n_2463), .B0 (n_6316), .B1(u3_rp_b3_b ), .Y (n_2565));
AOI22X1 g37602(.A0 (n_709), .A1 (n_2465), .B0 (n_6821), .B1(u6_rp_b3_b ), .Y (n_2566));
AOI22X1 g37601(.A0 (n_712), .A1 (n_3556), .B0 (n_145), .B1 (u4_rp_b3_b), .Y (n_3940));
AOI22X1 g37600(.A0 (n_639), .A1 (n_2468), .B0 (n_2567), .B1(u8_rp_b3_b ), .Y (n_2568));
AOI22X1 g37609(.A0 (in_slt_414), .A1 (n_4623), .B0 (in_slt_402), .B1(n_2368), .Y (n_5736));
NAND2X1 g37608(.A (n_2461), .B (n_2640), .Y (n_4630));
OAI21X1 g33777(.A0 (n_5044), .A1 (n_9100), .B0 (n_7750), .Y (n_9101));
OAI21X1 g33776(.A0 (n_5041), .A1 (n_9100), .B0 (n_7751), .Y (n_9102));
OAI21X1 g33812(.A0 (n_4903), .A1 (n_9034), .B0 (n_7716), .Y (n_9060));
OAI21X1 g33774(.A0 (n_4923), .A1 (n_9105), .B0 (n_7753), .Y (n_9104));
OAI21X1 g33773(.A0 (n_4924), .A1 (n_9105), .B0 (n_7754), .Y (n_9106));
OAI21X1 g33772(.A0 (n_4925), .A1 (n_9105), .B0 (n_7755), .Y (n_9107));
OAI21X1 g33770(.A0 (n_4926), .A1 (n_9110), .B0 (n_7757), .Y (n_9109));
OAI21X1 g33779(.A0 (n_5050), .A1 (n_9100), .B0 (n_7748), .Y (n_9098));
OAI21X1 g33778(.A0 (n_4922), .A1 (n_9100), .B0 (n_7749), .Y (n_9099));
NAND2X1 g38927(.A (u7_mem_b3_b_129 ), .B (n_1538), .Y (n_1529));
MX2X1 g38601(.A (u3_mem_b0_b_101 ), .B (wb_din_671), .S0 (n_3807), .Y(n_3811));
NAND2X1 g37463(.A (u13_ints_r_b8_b ), .B (n_3979), .Y (n_3970));
NAND2X1 g37462(.A (u13_ints_r_b7_b ), .B (n_3985), .Y (n_2579));
NAND2X1 g37461(.A (u13_ints_r_b6_b ), .B (n_3985), .Y (n_2580));
NAND2X1 g37460(.A (u13_ints_r_b5_b ), .B (n_3979), .Y (n_3971));
OAI21X1 g35875(.A0 (n_5563), .A1 (n_7115), .B0 (n_5880), .Y (n_6997));
NAND2X1 g37466(.A (n_5277), .B (crac_out_864), .Y (n_3968));
NAND2X1 g37465(.A (u13_ints_r_b25_b ), .B (n_4726), .Y (n_2613));
NAND2X1 g37464(.A (n_3979), .B (u13_ints_r_b9_b ), .Y (n_3969));
NAND2X1 g37469(.A (u13_ints_r_b12_b ), .B (n_3979), .Y (n_3966));
NAND2X1 g37468(.A (n_5277), .B (crac_out_863), .Y (n_3967));
CLKBUFX3 g41183(.A (n_1406), .Y (n_3935));
INVX1 g41184(.A (n_1899), .Y (n_4623));
INVX1 g41189(.A (n_1406), .Y (n_1899));
NAND2X1 g38925(.A (u7_mem_b3_b_124 ), .B (n_1538), .Y (n_1531));
AOI22X1 g37947(.A0 (n_5981), .A1 (n_940), .B0 (n_6005), .B1 (n_1316),.Y (n_3893));
NAND2X1 g38924(.A (u7_mem_b3_b ), .B (n_1538), .Y (n_1354));
INVX1 g42984(.A (n_1481), .Y (n_11059));
INVX1 g42633(.A (ic1_int_set_722), .Y (n_608));
INVX1 g42630(.A (u10_mem_b0_b_159 ), .Y (n_6386));
INVX1 g42631(.A (u9_mem_b3_b ), .Y (n_6924));
INVX1 g42636(.A (u11_mem_b3_b_64 ), .Y (n_6650));
INVX1 g42981(.A (n_1481), .Y (n_11069));
INVX1 g42634(.A (u9_mem_b1_b_120 ), .Y (n_6879));
MX2X1 g38761(.A (u3_mem_b0_b_96 ), .B (wb_din_666), .S0 (n_858), .Y(n_3574));
NAND2X1 g31601(.A (n_1715), .B (n_10054), .Y (n_10049));
NAND2X1 g31600(.A (n_2506), .B (n_10045), .Y (n_10050));
NAND2X1 g31603(.A (n_1863), .B (n_10010), .Y (n_10047));
NAND2X1 g31602(.A (n_2542), .B (n_10010), .Y (n_10048));
NAND2X1 g31605(.A (n_141), .B (n_10045), .Y (n_10044));
NAND2X1 g31604(.A (n_1766), .B (n_10045), .Y (n_10046));
NAND2X1 g31607(.A (n_35), .B (n_10054), .Y (n_10042));
NAND2X1 g31606(.A (n_1744), .B (n_10054), .Y (n_10043));
NAND2X1 g31609(.A (n_1561), .B (n_10045), .Y (n_10040));
NAND2X1 g31608(.A (n_198), .B (n_10045), .Y (n_10041));
OAI21X1 g35871(.A0 (n_5722), .A1 (n_11934), .B0 (n_6267), .Y(n_7046));
AND2X1 g41725(.A (u2_res_cnt_b0_b ), .B (u2_res_cnt_b2_b ), .Y (n_416));
NOR2X1 g41724(.A (u13_ints_r_b28_b ), .B (n_749), .Y (n_750));
NAND2X1 g41727(.A (wb_cyc_i), .B (wb_stb_i), .Y (n_2599));
INVX1 g41726(.A (n_2599), .Y (n_581));
INVX1 g35129(.A (n_7408), .Y (n_9290));
OAI21X1 g30958(.A0 (n_4752), .A1 (n_10450), .B0 (n_10066), .Y(n_10757));
OAI21X1 g30959(.A0 (n_5737), .A1 (n_10747), .B0 (n_10064), .Y(n_10756));
OAI21X1 g30956(.A0 (n_4762), .A1 (n_10450), .B0 (n_10069), .Y(n_10760));
OAI21X1 g30957(.A0 (n_4760), .A1 (n_10679), .B0 (n_10067), .Y(n_10758));
OAI21X1 g30954(.A0 (n_5378), .A1 (n_10450), .B0 (n_10072), .Y(n_10763));
OAI21X1 g30955(.A0 (n_5377), .A1 (n_10450), .B0 (n_10071), .Y(n_10762));
OAI21X1 g30952(.A0 (n_5740), .A1 (n_10747), .B0 (n_10075), .Y(n_10765));
OAI21X1 g30953(.A0 (n_5738), .A1 (n_10747), .B0 (n_10074), .Y(n_10764));
OAI21X1 g30950(.A0 (n_5379), .A1 (n_10679), .B0 (n_10078), .Y(n_10768));
OAI21X1 g30951(.A0 (n_5283), .A1 (n_10450), .B0 (n_10076), .Y(n_10766));
OAI21X1 g36730(.A0 (n_2513), .A1 (u11_wp_b1_b ), .B0 (n_1816), .Y(n_4073));
MX2X1 g36731(.A (u10_mem_b0_b_167 ), .B (n_5418), .S0 (n_6341), .Y(n_5419));
MX2X1 g36732(.A (u11_mem_b0_b_168 ), .B (n_5410), .S0 (n_6359), .Y(n_5416));
MX2X1 g36733(.A (u10_mem_b0_b_168 ), .B (n_5422), .S0 (n_6341), .Y(n_5415));
XOR2X1 g36734(.A (u26_ps_cnt_b5_b ), .B (n_1775), .Y (n_4827));
MX2X1 g36735(.A (u11_mem_b1_b_136 ), .B (n_5413), .S0 (n_5405), .Y(n_5414));
MX2X1 g36737(.A (u11_mem_b2_b_105 ), .B (n_5413), .S0 (n_5409), .Y(n_5412));
MX2X1 g36738(.A (u11_mem_b2_b_106 ), .B (n_5410), .S0 (n_5409), .Y(n_5411));
MX2X1 g36739(.A (u9_mem_b1_b_137 ), .B (n_5733), .S0 (n_5730), .Y(n_5731));
NAND2X1 g38844(.A (u5_mem_b3_b_144 ), .B (n_3543), .Y (n_2444));
INVX1 g42186(.A (u26_cnt_b1_b ), .Y (n_37));
INVX1 g42180(.A (u9_mem_b0_b_163 ), .Y (n_6398));
INVX1 g42181(.A (u11_mem_b3_b_77 ), .Y (n_5526));
INVX1 g42182(.A (u10_mem_b2_b_111 ), .Y (n_9));
INVX4 g41686(.A (n_1364), .Y (n_3339));
INVX1 g39609(.A (n_4776), .Y (n_3060));
NAND2X1 g38845(.A (u5_mem_b3_b_130 ), .B (n_1543), .Y (n_1326));
NOR2X1 g39603(.A (n_3089), .B (n_2782), .Y (n_3067));
INVX1 g35384(.A (i6_status_1042), .Y (n_7030));
NAND2X1 g39604(.A (n_11789), .B (u8_mem_b0_b_121 ), .Y (n_3066));
INVX1 g39607(.A (n_4759), .Y (n_3061));
INVX1 g35387(.A (i4_status_1032), .Y (n_6720));
MX2X1 g34910(.A (i4_full), .B (u14_u7_full_empty_r), .S0 (n_7357), .Y(n_7557));
MX2X1 g38765(.A (u8_mem_b0_b_97 ), .B (wb_din_667), .S0 (n_3826), .Y(n_3570));
NAND2X1 g38846(.A (u5_mem_b3_b_132 ), .B (n_1543), .Y (n_1542));
MX2X1 g34911(.A (i6_full), .B (u14_u8_full_empty_r), .S0 (n_7388), .Y(n_8213));
NAND2X1 g38847(.A (u5_mem_b3_b_145 ), .B (n_3543), .Y (n_3545));
NAND2X1 g39889(.A (n_11798), .B (u8_mem_b0_b ), .Y (n_11467));
NAND2X1 g34659(.A (u6_mem_b2_b_32 ), .B (n_7758), .Y (n_7766));
NAND2X1 g34658(.A (u6_mem_b2_b_31 ), .B (n_7758), .Y (n_7767));
NAND2X1 g34655(.A (u6_mem_b2_b_30 ), .B (n_7758), .Y (n_7770));
OAI21X1 g33974(.A0 (n_4483), .A1 (n_8933), .B0 (n_8062), .Y (n_8849));
MX2X1 g33977(.A (u3_mem_b0_b_112 ), .B (n_3834), .S0 (n_8700), .Y(n_8842));
OAI21X1 g33976(.A0 (n_4487), .A1 (n_8933), .B0 (n_8067), .Y (n_8845));
OAI21X1 g33971(.A0 (n_4856), .A1 (n_8856), .B0 (n_7562), .Y (n_8852));
OAI21X1 g33970(.A0 (n_4477), .A1 (n_8868), .B0 (n_7563), .Y (n_8854));
NAND2X1 g34653(.A (u6_mem_b2_b_56 ), .B (n_7758), .Y (n_7772));
NAND2X1 g34652(.A (u6_mem_b2_b_55 ), .B (n_7758), .Y (n_7773));
NAND2X1 g34556(.A (u5_mem_b3_b_131 ), .B (n_7870), .Y (n_7871));
INVX2 g41041(.A (n_821), .Y (n_1027));
NAND2X1 g39584(.A (n_2344), .B (in_slt_428), .Y (n_2280));
NAND2X1 g34557(.A (u5_mem_b3_b_132 ), .B (n_7870), .Y (n_7869));
NAND2X1 g34554(.A (u5_mem_b2_b_37 ), .B (n_7870), .Y (n_7873));
NAND3X1 g45468(.A (n_11924), .B (n_11658), .C (n_4251), .Y (n_11925));
NAND2X1 g34555(.A (u5_mem_b3_b ), .B (n_7870), .Y (n_7872));
NAND2X1 g34552(.A (u5_mem_b2_b_35 ), .B (n_7870), .Y (n_7875));
NAND2X1 g38841(.A (u4_mem_b3_b_133 ), .B (n_3546), .Y (n_3547));
NAND2X1 g34553(.A (u5_mem_b2_b_36 ), .B (n_7870), .Y (n_7874));
NAND2X1 g34387(.A (u4_mem_b2_b_38 ), .B (n_7984), .Y (n_8017));
NAND2X1 g34386(.A (u4_mem_b2_b ), .B (n_7984), .Y (n_8018));
NAND2X1 g34385(.A (n_6683), .B (n_7463), .Y (n_8229));
NAND2X1 g34384(.A (u4_mem_b1_b_68 ), .B (n_7984), .Y (n_8019));
NAND2X1 g34383(.A (u4_mem_b1_b_67 ), .B (n_7984), .Y (n_8020));
NAND2X1 g34550(.A (u5_mem_b2_b_33 ), .B (n_7870), .Y (n_7877));
NAND2X1 g34381(.A (u4_mem_b1_b_65 ), .B (n_7984), .Y (n_8022));
NAND2X1 g34380(.A (u4_mem_b1_b_64 ), .B (n_7984), .Y (n_8023));
NAND2X1 g34551(.A (u5_mem_b2_b_34 ), .B (n_7870), .Y (n_7876));
NAND2X1 g34389(.A (u4_mem_b2_b_40 ), .B (n_7984), .Y (n_8015));
NAND2X1 g34388(.A (u4_mem_b2_b_39 ), .B (n_7984), .Y (n_8016));
NAND2X1 g34478(.A (u3_mem_b2_b_49 ), .B (n_8101), .Y (n_7946));
MX2X1 g38769(.A (u7_mem_b0_b_91 ), .B (wb_din_661), .S0 (n_913), .Y(n_3566));
NAND2X1 g34471(.A (u4_mem_b3_b_130 ), .B (n_7984), .Y (n_7950));
NAND2X1 g34470(.A (u4_mem_b3_b_129 ), .B (n_7984), .Y (n_7951));
NOR2X1 g34473(.A (n_1419), .B (n_7984), .Y (n_8227));
NAND2X1 g34472(.A (u8_mem_b1_b_82 ), .B (n_7976), .Y (n_7949));
INVX4 g34475(.A (n_7445), .Y (n_8519));
NAND2X1 g34474(.A (u8_mem_b1_b_71 ), .B (n_7976), .Y (n_7948));
NAND2X1 g34477(.A (u3_mem_b1_b_79 ), .B (n_8101), .Y (n_7947));
NAND2X1 g34476(.A (n_7444), .B (n_6044), .Y (n_7445));
MX2X1 g34009(.A (u4_mem_b0_b_96 ), .B (n_3755), .S0 (n_7499), .Y(n_8812));
AOI22X1 g37652(.A0 (n_6628), .A1 (n_1835), .B0 (n_6559), .B1(n_1760), .Y (n_1707));
NAND2X1 g38843(.A (u5_mem_b3_b_129 ), .B (n_1543), .Y (n_1544));
OAI21X1 g45872(.A0 (n_12605), .A1 (n_12606), .B0 (n_12609), .Y(n_12610));
INVX1 g42099(.A (u10_mem_b0_b_170 ), .Y (n_1244));
MX2X1 g38642(.A (u8_mem_b0_b_120 ), .B (wb_din_690), .S0 (n_3826), .Y(n_3748));
AOI21X1 g38215(.A0 (u4_mem_b3_b_150 ), .A1 (n_5106), .B0 (n_3506), .Y(n_5080));
NAND2X1 g39585(.A (n_2325), .B (in_slt_451), .Y (n_2279));
MX2X1 g38643(.A (u8_mem_b0_b_92 ), .B (wb_din_662), .S0 (n_3826), .Y(n_3746));
NOR2X1 g39283(.A (u10_mem_b1_b_140 ), .B (n_2364), .Y (n_2332));
NAND2X1 g32734(.A (n_348), .B (n_10605), .Y (n_12063));
NAND2X1 g32735(.A (n_297), .B (n_10583), .Y (n_11628));
NAND2X1 g32736(.A (n_200), .B (n_10605), .Y (n_11995));
NAND2X1 g32737(.A (n_208), .B (n_10583), .Y (n_11622));
AOI21X1 g32730(.A0 (n_6185), .A1 (n_6151), .B0 (n_10605), .Y(n_10589));
NAND2X1 g32731(.A (n_203), .B (n_10583), .Y (n_11618));
AOI21X1 g32732(.A0 (n_6179), .A1 (n_6177), .B0 (n_10605), .Y(n_10587));
NAND2X1 g32733(.A (n_263), .B (n_10583), .Y (n_11620));
MX2X1 g38640(.A (u3_mem_b0_b_99 ), .B (wb_din_669), .S0 (n_858), .Y(n_3751));
NAND2X1 g32738(.A (n_150), .B (n_10583), .Y (n_11624));
NAND2X1 g32739(.A (n_211), .B (n_10605), .Y (n_11732));
NAND2X1 g36650(.A (n_5258), .B (n_3970), .Y (n_5780));
INVX1 g43067(.A (u6_wp_b0_b ), .Y (n_706));
AOI21X1 g38408(.A0 (u6_mem_b1_b_76 ), .A1 (n_5112), .B0 (n_2737), .Y(n_4945));
AOI21X1 g38409(.A0 (u6_mem_b1_b_75 ), .A1 (n_5112), .B0 (n_2787), .Y(n_4944));
AOI21X1 g38159(.A0 (u4_mem_b2_b_50 ), .A1 (n_4439), .B0 (n_1991), .Y(n_4427));
AOI21X1 g38157(.A0 (u6_mem_b1_b_67 ), .A1 (n_5019), .B0 (n_2657), .Y(n_5111));
AOI21X1 g38154(.A0 (u4_mem_b2_b_46 ), .A1 (n_4439), .B0 (n_2102), .Y(n_4431));
AOI21X1 g38407(.A0 (u6_mem_b1_b_72 ), .A1 (n_5019), .B0 (n_2682), .Y(n_4946));
AOI21X1 g38152(.A0 (u4_mem_b2_b_45 ), .A1 (n_4439), .B0 (n_1976), .Y(n_4432));
AOI21X1 g38153(.A0 (u6_mem_b1_b_66 ), .A1 (n_5112), .B0 (n_2690), .Y(n_5113));
AOI21X1 g38150(.A0 (u4_mem_b2_b_44 ), .A1 (n_4439), .B0 (n_2110), .Y(n_4433));
AOI21X1 g38151(.A0 (u4_mem_b3_b ), .A1 (n_5106), .B0 (n_3313), .Y(n_5114));
MX2X1 g31343(.A (n_6334), .B (n_6333), .S0 (n_10137), .Y (n_10120));
NAND2X1 g38848(.A (u7_mem_b3_b_147 ), .B (n_1546), .Y (n_1328));
MX2X1 g38646(.A (u5_mem_b0_b_100 ), .B (wb_din_670), .S0 (n_3720), .Y(n_3739));
NAND2X1 g38970(.A (u3_mem_b3_b_123 ), .B (n_1517), .Y (n_1378));
NOR2X1 g40118(.A (n_2470), .B (n_2801), .Y (n_2116));
MX2X1 g31344(.A (n_5946), .B (n_5945), .S0 (n_10137), .Y (n_10119));
NAND2X1 g38971(.A (u8_mem_b3_b_134 ), .B (n_2468), .Y (n_2390));
NOR2X1 g40115(.A (n_2681), .B (n_2118), .Y (n_2119));
NOR2X1 g40114(.A (n_2120), .B (n_2790), .Y (n_2121));
NOR2X1 g40117(.A (n_2103), .B (n_2735), .Y (n_2117));
NOR2X1 g40116(.A (n_2784), .B (n_2765), .Y (n_2758));
NOR2X1 g40111(.A (n_2470), .B (n_2748), .Y (n_2123));
AOI21X1 g37252(.A0 (n_5352), .A1 (n_6594), .B0 (n_3956), .Y (n_5353));
NOR2X1 g40113(.A (n_2818), .B (n_2118), .Y (n_2122));
NOR2X1 g40112(.A (n_2759), .B (n_2691), .Y (n_2760));
NAND2X1 g38973(.A (u6_mem_b3_b_148 ), .B (n_2465), .Y (n_2388));
MX2X1 g38647(.A (u5_mem_b0_b_101 ), .B (wb_din_671), .S0 (n_3720), .Y(n_3737));
NAND2X1 g38974(.A (u8_mem_b3_b_136 ), .B (n_2468), .Y (n_2387));
AOI21X1 g37255(.A0 (n_5506), .A1 (n_6594), .B0 (n_4656), .Y (n_5507));
AOI21X1 g37708(.A0 (n_6007), .A1 (n_1316), .B0 (n_2336), .Y (n_3923));
NAND2X1 g37709(.A (n_3550), .B (n_3328), .Y (n_4603));
AOI22X1 g37706(.A0 (in_slt3), .A1 (n_1406), .B0 (u9_din_tmp1), .B1(n_2368), .Y (n_4605));
MX2X1 g38644(.A (u3_mem_b0_b_93 ), .B (wb_din_663), .S0 (n_3807), .Y(n_3744));
NAND2X1 g38979(.A (u8_mem_b3_b_123 ), .B (n_2468), .Y (n_2384));
NAND2X1 g36383(.A (n_5895), .B (n_2567), .Y (n_5913));
MX2X1 g38645(.A (u5_mem_b0_b ), .B (wb_din), .S0 (n_3720), .Y(n_3741));
NAND2X1 g39829(.A (u4_mem_b1_b ), .B (n_12252), .Y (n_11671));
AOI22X1 g37701(.A0 (u10_din_tmp_46), .A1 (n_3339), .B0 (n_3911), .B1(in_slt_425), .Y (n_3928));
NAND2X1 g39533(.A (n_2344), .B (in_slt_420), .Y (n_2290));
NOR2X1 g39532(.A (n_3117), .B (n_2712), .Y (n_3111));
OAI21X1 g45464(.A0 (n_11922), .A1 (n_11928), .B0 (n_12149), .Y(n_12006));
NAND2X1 g39531(.A (u7_mem_b2_b_42 ), .B (n_12645), .Y (n_3112));
AOI22X1 g37818(.A0 (n_277), .A1 (n_1575), .B0 (n_5490), .B1 (n_1831),.Y (n_1617));
AOI21X1 g30847(.A0 (n_10625), .A1 (n_10207), .B0 (n_5825), .Y(n_11074));
AOI22X1 g37812(.A0 (n_6406), .A1 (n_2530), .B0 (n_6607), .B1(n_2544), .Y (n_2528));
NAND2X1 g37813(.A (n_1536), .B (n_4121), .Y (n_5210));
NAND2X1 g37810(.A (n_4198), .B (n_3173), .Y (n_5211));
AOI22X1 g37811(.A0 (n_339), .A1 (n_1643), .B0 (n_5526), .B1 (n_1831),.Y (n_1625));
AOI22X1 g37816(.A0 (n_2558), .A1 (n_6333), .B0 (n_6562), .B1(n_1316), .Y (n_1235));
AOI22X1 g37817(.A0 (n_1756), .A1 (n_1620), .B0 (n_1619), .B1(n_1643), .Y (n_1621));
AOI22X1 g37814(.A0 (n_279), .A1 (n_1575), .B0 (n_5488), .B1 (n_1831),.Y (n_1623));
NAND2X1 g39536(.A (u3_mem_b1_b_87 ), .B (n_3316), .Y (n_3107));
INVX2 g41538(.A (n_9719), .Y (n_7256));
MX2X1 g33128(.A (ic2_cfg_1050), .B (wb_din_683), .S0 (n_8611), .Y(n_8589));
NAND2X1 g39535(.A (n_12839), .B (u4_mem_b0_b_91 ), .Y (n_3108));
AOI21X1 g45465(.A0 (n_6322), .A1 (n_6124), .B0 (n_7324), .Y(n_11922));
MX2X1 g33122(.A (n_4683), .B (wb_din_678), .S0 (n_8611), .Y (n_8604));
MX2X1 g33123(.A (n_4706), .B (wb_din_679), .S0 (n_8611), .Y (n_8601));
MX2X1 g33120(.A (n_11772), .B (wb_din_676), .S0 (n_8611), .Y(n_8608));
MX2X1 g33121(.A (ic2_cfg_1044), .B (wb_din_677), .S0 (n_8611), .Y(n_8606));
MX2X1 g33126(.A (n_5588), .B (wb_din_681), .S0 (n_8611), .Y (n_8594));
MX2X1 g33127(.A (ic2_cfg_1049), .B (wb_din_682), .S0 (n_8611), .Y(n_8592));
MX2X1 g33124(.A (ic0_cfg_1024), .B (wb_din_661), .S0 (n_8611), .Y(n_8599));
MX2X1 g33125(.A (n_5788), .B (wb_din_680), .S0 (n_8611), .Y (n_8597));
MX2X1 g31142(.A (n_6613), .B (n_6612), .S0 (n_9724), .Y (n_10649));
MX2X1 g31143(.A (n_6583), .B (n_6581), .S0 (n_10747), .Y (n_10254));
MX2X1 g31140(.A (n_6451), .B (n_6450), .S0 (n_10235), .Y (n_10258));
MX2X1 g31141(.A (n_6506), .B (n_6505), .S0 (n_10747), .Y (n_10256));
MX2X1 g31146(.A (n_6921), .B (n_6919), .S0 (n_10250), .Y (n_10251));
MX2X1 g31147(.A (n_6608), .B (n_6607), .S0 (n_10315), .Y (n_10249));
MX2X1 g31144(.A (n_6923), .B (n_6922), .S0 (n_10235), .Y (n_10253));
MX2X1 g31145(.A (n_6953), .B (n_6951), .S0 (n_10235), .Y (n_10252));
MX2X1 g31148(.A (n_6917), .B (n_6915), .S0 (n_10250), .Y (n_10247));
MX2X1 g31149(.A (n_6892), .B (n_6890), .S0 (n_10277), .Y (n_10245));
INVX1 g39647(.A (n_5284), .Y (n_4153));
NAND2X1 g39317(.A (u3_mem_b1_b_66 ), .B (n_3316), .Y (n_3278));
NOR2X1 g39316(.A (n_5102), .B (n_2748), .Y (n_3279));
AOI21X1 g38574(.A0 (u3_mem_b1_b_82 ), .A1 (n_5148), .B0 (n_2822), .Y(n_4858));
NAND2X1 g39858(.A (in_slt_408), .B (n_2368), .Y (n_4753));
NOR2X1 g39315(.A (n_3486), .B (n_2804), .Y (n_3280));
NAND2X1 g39854(.A (u8_mem_b2_b_43 ), .B (n_2362), .Y (n_2237));
MX2X1 g38649(.A (u5_mem_b0_b_104 ), .B (wb_din_674), .S0 (n_3720), .Y(n_3734));
NAND2X1 g39856(.A (u8_mem_b2_b_30 ), .B (n_2366), .Y (n_11501));
NAND2X1 g39314(.A (u8_mem_b1_b_80 ), .B (n_12291), .Y (n_3282));
NAND2X1 g39850(.A (u3_mem_b1_b_82 ), .B (n_3316), .Y (n_2923));
AOI21X1 g38576(.A0 (u3_mem_b1_b_83 ), .A1 (n_5157), .B0 (n_2663), .Y(n_4857));
NOR2X1 g39853(.A (n_2755), .B (n_1488), .Y (n_1464));
OAI21X1 g37381(.A0 (u9_mem_b0_b_170 ), .A1 (n_6856), .B0 (n_4673), .Y(n_5484));
INVX1 g42329(.A (n_12331), .Y (n_1921));
INVX1 g41921(.A (u2_to_cnt_b3_b ), .Y (n_703));
AOI21X1 g38571(.A0 (u3_mem_b1_b_79 ), .A1 (n_5148), .B0 (n_2815), .Y(n_4861));
OAI21X1 g37384(.A0 (u9_mem_b0_b_174 ), .A1 (n_5480), .B0 (n_4659), .Y(n_5481));
NAND2X1 g39649(.A (n_12389), .B (u4_mem_b0_b_121 ), .Y (n_3036));
OAI21X1 g33584(.A0 (n_5089), .A1 (n_8318), .B0 (n_7969), .Y (n_9342));
AOI21X1 g38573(.A0 (u3_mem_b3_b ), .A1 (n_5138), .B0 (n_2937), .Y(n_4859));
NAND2X1 g38814(.A (u7_mem_b3_b_123 ), .B (n_1538), .Y (n_1275));
INVX1 g41925(.A (u10_mem_b0_b_155 ), .Y (n_6331));
INVX1 g41924(.A (u9_mem_b3_b_60 ), .Y (n_6895));
NAND4X1 g36920(.A (n_11443), .B (n_1319), .C (n_11444), .D (n_1335),.Y (n_5869));
INVX1 g36924(.A (n_5707), .Y (n_5708));
AOI22X1 g35713(.A0 (n_6686), .A1 (i6_dout_650), .B0 (i4_dout_619),.B1 (n_7297), .Y (n_7012));
AOI22X1 g35712(.A0 (n_6686), .A1 (i6_dout_649), .B0 (i4_dout_618),.B1 (n_7297), .Y (n_6673));
AOI22X1 g35711(.A0 (n_6686), .A1 (i6_dout_645), .B0 (i4_dout_614),.B1 (n_7297), .Y (n_7112));
XOR2X1 g35717(.A (n_5442), .B (n_4072), .Y (n_5638));
AOI21X1 g35716(.A0 (i4_dout_625), .A1 (n_7468), .B0 (n_7111), .Y(n_7302));
AOI21X1 g35715(.A0 (i4_dout_624), .A1 (n_7297), .B0 (n_7151), .Y(n_7298));
AOI21X1 g35714(.A0 (i4_dout_623), .A1 (n_7468), .B0 (n_7107), .Y(n_7296));
XOR2X1 g35719(.A (n_2612), .B (n_4104), .Y (n_5431));
XOR2X1 g35718(.A (n_4851), .B (n_2611), .Y (n_5449));
INVX1 g35248(.A (o3_status_962), .Y (n_7037));
INVX1 g42370(.A (u10_mem_b1_b_147 ), .Y (n_2538));
INVX1 g42377(.A (u11_mem_b1_b_139 ), .Y (n_339));
INVX1 g42375(.A (u9_mem_b2_b_90 ), .Y (n_6888));
CLKBUFX1 g40936(.A (n_931), .Y (n_5424));
INVX4 g46004(.A (n_12735), .Y (n_12825));
INVX1 g42379(.A (n_9833), .Y (n_10916));
INVX1 g43022(.A (u9_mem_b2_b_99 ), .Y (n_6495));
INVX2 g32948(.A (n_9720), .Y (n_10385));
INVX1 g43024(.A (u11_mem_b2_b_106 ), .Y (n_288));
INVX1 g43026(.A (u9_mem_b2_b_104 ), .Y (n_6935));
INVX2 g43028(.A (n_1875), .Y (n_11086));
INVX4 g32942(.A (n_9905), .Y (n_10880));
INVX4 g32947(.A (n_9720), .Y (n_10376));
NAND2X1 g39795(.A (u4_mem_b2_b_44 ), .B (n_12087), .Y (n_2246));
INVX4 g32945(.A (n_9720), .Y (n_9818));
INVX2 g32944(.A (n_9818), .Y (n_9905));
NAND2X1 g39149(.A (in_slt_402), .B (n_3415), .Y (n_3416));
NOR2X1 g40289(.A (n_2702), .B (n_1985), .Y (n_1986));
NOR2X1 g40288(.A (n_3008), .B (n_2067), .Y (n_1987));
NAND2X1 g39142(.A (n_12389), .B (u4_mem_b0_b_119 ), .Y (n_3422));
INVX1 g39143(.A (n_4749), .Y (n_3420));
NOR2X1 g39140(.A (n_3089), .B (n_2707), .Y (n_3425));
NAND2X1 g39141(.A (u6_mem_b2_b_54 ), .B (n_3423), .Y (n_3424));
NAND2X1 g39146(.A (u7_mem_b1_b_76 ), .B (n_4225), .Y (n_4226));
NAND2X1 g39147(.A (u6_mem_b1_b_84 ), .B (n_4253), .Y (n_4224));
NOR2X1 g40283(.A (n_1147), .B (n_2681), .Y (n_2682));
NAND2X1 g39145(.A (u8_mem_b1_b_82 ), .B (n_12291), .Y (n_3419));
MX2X1 g34040(.A (u5_mem_b0_b_94 ), .B (n_3696), .S0 (n_7496), .Y(n_9420));
MX2X1 g34041(.A (u5_mem_b0_b_95 ), .B (n_3690), .S0 (n_7496), .Y(n_8784));
MX2X1 g34042(.A (u5_mem_b0_b_96 ), .B (n_3688), .S0 (n_7496), .Y(n_8783));
MX2X1 g34043(.A (u5_mem_b0_b_97 ), .B (n_3694), .S0 (n_7496), .Y(n_9419));
MX2X1 g34044(.A (u5_mem_b0_b_98 ), .B (n_3693), .S0 (n_7496), .Y(n_8782));
MX2X1 g34045(.A (u5_mem_b0_b_99 ), .B (n_3692), .S0 (n_7496), .Y(n_9417));
MX2X1 g34046(.A (u3_mem_b0_b_92 ), .B (n_3820), .S0 (n_8700), .Y(n_9416));
MX2X1 g34047(.A (u6_mem_b0_b ), .B (n_3683), .S0 (n_7505), .Y(n_8781));
MX2X1 g34048(.A (u6_mem_b0_b_100 ), .B (n_3682), .S0 (n_7505), .Y(n_8780));
MX2X1 g34049(.A (u6_mem_b0_b_101 ), .B (n_3565), .S0 (n_7505), .Y(n_8779));
AOI21X1 g40388(.A0 (u5_rp_b3_b ), .A1 (u5_wp_b2_b ), .B0 (n_412), .Y(n_968));
INVX4 g46005(.A (n_12244), .Y (n_12839));
NAND2X1 g39884(.A (u7_mem_b2_b_36 ), .B (n_12645), .Y (n_3848));
AOI21X1 g38325(.A0 (u6_mem_b2_b_57 ), .A1 (n_4544), .B0 (n_1953), .Y(n_4358));
AOI21X1 g40389(.A0 (u9_rp_b0_b ), .A1 (n_4074), .B0 (n_1054), .Y(n_4851));
NAND2X1 g29930(.A (n_11123), .B (u16_u4_dma_req_r1), .Y (n_11171));
NAND2X1 g29931(.A (n_11122), .B (u16_u5_dma_req_r1), .Y (n_11170));
AOI21X1 g38365(.A0 (u5_mem_b3_b_152 ), .A1 (n_5000), .B0 (n_3118), .Y(n_4972));
AOI21X1 g38364(.A0 (u6_mem_b1_b_78 ), .A1 (n_5019), .B0 (n_2821), .Y(n_4973));
AOI21X1 g38367(.A0 (u5_mem_b3_b_125 ), .A1 (n_5000), .B0 (n_3114), .Y(n_4970));
AOI21X1 g38366(.A0 (u5_mem_b3_b_124 ), .A1 (n_5000), .B0 (n_3116), .Y(n_4971));
AOI21X1 g38361(.A0 (u5_mem_b3_b_123 ), .A1 (n_4996), .B0 (n_3353), .Y(n_4976));
AOI21X1 g38360(.A0 (u5_mem_b3_b_150 ), .A1 (n_5000), .B0 (n_3010), .Y(n_4977));
AOI21X1 g38363(.A0 (u5_mem_b3_b_151 ), .A1 (n_5000), .B0 (n_3018), .Y(n_4974));
AOI21X1 g38362(.A0 (u7_mem_b1_b_83 ), .A1 (n_5118), .B0 (n_2791), .Y(n_4975));
AOI22X1 g37669(.A0 (n_2502), .A1 (n_1701), .B0 (n_1700), .B1(n_1835), .Y (n_1702));
AOI22X1 g37668(.A0 (in_slt_400), .A1 (n_1406), .B0 (u9_din_tmp_45),.B1 (n_4616), .Y (n_4617));
AOI21X1 g38369(.A0 (u5_mem_b3_b_128 ), .A1 (n_4996), .B0 (n_3111), .Y(n_4968));
AOI21X1 g38368(.A0 (u5_mem_b3_b_126 ), .A1 (n_5000), .B0 (n_3027), .Y(n_4969));
OAI21X1 g33711(.A0 (n_4944), .A1 (n_9182), .B0 (n_7823), .Y (n_9183));
OAI21X1 g33710(.A0 (n_4941), .A1 (n_9161), .B0 (n_7824), .Y (n_9185));
OAI21X1 g33713(.A0 (n_4967), .A1 (n_9182), .B0 (n_7821), .Y (n_9179));
OAI21X1 g33712(.A0 (n_4945), .A1 (n_9182), .B0 (n_7822), .Y (n_9181));
OAI21X1 g33715(.A0 (n_4943), .A1 (n_9161), .B0 (n_7817), .Y (n_9176));
OAI21X1 g33714(.A0 (n_4973), .A1 (n_9182), .B0 (n_7819), .Y (n_9177));
OAI21X1 g33717(.A0 (n_5003), .A1 (n_9139), .B0 (n_7813), .Y (n_9174));
OAI21X1 g33716(.A0 (n_4942), .A1 (n_9110), .B0 (n_7815), .Y (n_9175));
OAI21X1 g33719(.A0 (n_5007), .A1 (n_9170), .B0 (n_7811), .Y (n_9172));
OAI21X1 g33718(.A0 (n_5004), .A1 (n_9161), .B0 (n_7812), .Y (n_9173));
NAND2X1 g37489(.A (n_5480), .B (n_3363), .Y (n_4670));
NAND2X1 g37488(.A (n_5480), .B (n_3420), .Y (n_4671));
NAND2X1 g37485(.A (n_1262), .B (n_1006), .Y (n_1263));
NOR2X1 g37484(.A (n_5317), .B (n_6649), .Y (n_4675));
NAND2X1 g37487(.A (n_5480), .B (n_3470), .Y (n_4672));
NAND2X1 g37486(.A (n_5480), .B (n_2895), .Y (n_4673));
INVX1 g37481(.A (n_2576), .Y (n_4676));
CLKBUFX3 g37480(.A (n_4676), .Y (n_6700));
NAND2X1 g37483(.A (n_5656), .B (n_4232), .Y (n_5246));
NAND2X1 g37482(.A (n_2575), .B (n_2574), .Y (n_2576));
CLKBUFX1 g46006(.A (n_12846), .Y (n_12845));
NOR2X1 g36538(.A (i3_status), .B (n_11563), .Y (n_5595));
NAND2X1 g36539(.A (n_6211), .B (n_6773), .Y (n_6212));
NOR2X1 g36536(.A (o9_status), .B (n_12585), .Y (n_5436));
NAND2X1 g36537(.A (n_12481), .B (n_6773), .Y (n_6215));
NAND2X1 g36534(.A (n_6186), .B (n_634), .Y (n_6218));
NAND2X1 g36535(.A (n_6216), .B (n_6773), .Y (n_6217));
NOR2X1 g36532(.A (o8_status), .B (n_5825), .Y (n_5826));
NAND2X1 g36533(.A (n_5823), .B (n_6259), .Y (n_5824));
NAND2X1 g36530(.A (n_12531), .B (n_6777), .Y (n_6778));
NOR2X1 g36531(.A (o7_status), .B (n_5827), .Y (n_5828));
INVX1 g42618(.A (u9_mem_b2_b_96 ), .Y (n_6893));
INVX1 g42969(.A (u11_mem_b1_b_119 ), .Y (n_6500));
INVX1 g42966(.A (u26_ps_cnt_b0_b ), .Y (n_529));
INVX1 g42962(.A (u6_wp_b1_b ), .Y (n_751));
INVX1 g42960(.A (n_751), .Y (n_7048));
NAND2X1 g31629(.A (n_5350), .B (n_10019), .Y (n_10014));
NAND2X1 g31628(.A (n_5365), .B (n_10019), .Y (n_10015));
NAND2X1 g31623(.A (n_5333), .B (n_10019), .Y (n_10022));
NAND2X1 g31622(.A (n_5372), .B (n_10019), .Y (n_10023));
NAND2X1 g31621(.A (n_5343), .B (n_10024), .Y (n_10025));
NAND2X1 g31620(.A (n_5374), .B (n_10019), .Y (n_10026));
NAND2X1 g31627(.A (n_5345), .B (n_10024), .Y (n_10016));
NAND2X1 g31626(.A (n_5347), .B (n_10024), .Y (n_10017));
NAND2X1 g31625(.A (n_5367), .B (n_10019), .Y (n_10018));
NAND2X1 g31624(.A (n_5302), .B (n_10019), .Y (n_10020));
OAI21X1 g30978(.A0 (n_4779), .A1 (n_10738), .B0 (n_10043), .Y(n_10730));
OAI21X1 g30979(.A0 (n_4748), .A1 (n_10738), .B0 (n_10042), .Y(n_10728));
NOR2X1 g41709(.A (wb_we_i), .B (u12_re2), .Y (n_1006));
AOI22X1 g35700(.A0 (n_6686), .A1 (i6_dout_632), .B0 (i3_dout_570),.B1 (n_6700), .Y (n_6684));
OAI21X1 g30970(.A0 (n_4785), .A1 (n_10738), .B0 (n_10053), .Y(n_10742));
OAI21X1 g30971(.A0 (n_4784), .A1 (n_10747), .B0 (n_10052), .Y(n_10740));
OAI21X1 g30972(.A0 (n_4782), .A1 (n_10738), .B0 (n_10050), .Y(n_10739));
OAI21X1 g30973(.A0 (n_4781), .A1 (n_10747), .B0 (n_10049), .Y(n_10737));
OAI21X1 g30974(.A0 (n_5331), .A1 (n_10450), .B0 (n_10048), .Y(n_10735));
OAI21X1 g30975(.A0 (n_5340), .A1 (n_10679), .B0 (n_10047), .Y(n_10733));
OAI21X1 g30976(.A0 (n_5735), .A1 (n_10019), .B0 (n_10046), .Y(n_10732));
OAI21X1 g30977(.A0 (n_5734), .A1 (n_10747), .B0 (n_10044), .Y(n_10731));
XOR2X1 g36750(.A (u2_to_cnt_b0_b ), .B (n_5630), .Y (n_5403));
INVX1 g36757(.A (o7_status), .Y (n_5400));
INVX1 g45390(.A (ic1_cfg), .Y (n_11612));
OAI21X1 g33838(.A0 (n_5045), .A1 (n_9022), .B0 (n_8089), .Y (n_9023));
MX2X1 g31089(.A (n_6667), .B (n_6666), .S0 (n_10137), .Y (n_10322));
MX2X1 g31088(.A (n_6669), .B (n_6668), .S0 (n_10137), .Y (n_10323));
MX2X1 g31087(.A (n_6611), .B (n_6610), .S0 (n_10137), .Y (n_10325));
MX2X1 g31086(.A (n_6036), .B (n_6035), .S0 (n_10537), .Y (n_10654));
MX2X1 g31085(.A (n_5999), .B (n_5998), .S0 (n_10137), .Y (n_10326));
MX2X1 g31084(.A (n_6651), .B (n_6650), .S0 (n_10537), .Y (n_10655));
AOI21X1 g31083(.A0 (n_11889), .A1 (u7_rp_b3_b ), .B0 (n_9967), .Y(n_10657));
AOI21X1 g31082(.A0 (n_11891), .A1 (u6_rp_b3_b ), .B0 (n_9969), .Y(n_10659));
MX2X1 g31081(.A (u5_rp_b3_b ), .B (n_4645), .S0 (n_10327), .Y(n_10328));
MX2X1 g31080(.A (u4_rp_b3_b ), .B (n_5467), .S0 (n_10329), .Y(n_10330));
NAND2X1 g39447(.A (u5_mem_b1_b_83 ), .B (n_3239), .Y (n_3176));
NAND2X1 g39446(.A (u7_mem_b1_b_67 ), .B (n_4130), .Y (n_4190));
NAND2X1 g39445(.A (u7_mem_b1_b_81 ), .B (n_4130), .Y (n_4191));
NOR2X1 g39444(.A (n_5059), .B (n_2732), .Y (n_3177));
NOR2X1 g39443(.A (n_5059), .B (n_2831), .Y (n_3180));
NAND2X1 g39442(.A (u3_mem_b1_b_75 ), .B (n_3316), .Y (n_3181));
OR2X1 g39441(.A (n_12604), .B (n_3559), .Y (n_2298));
NAND2X1 g39440(.A (u8_mem_b2_b_39 ), .B (n_2362), .Y (n_2299));
NAND2X1 g39449(.A (n_3252), .B (u7_mem_b0_b_117 ), .Y (n_3173));
NOR2X1 g39448(.A (n_3332), .B (n_2790), .Y (n_3175));
NAND2X1 g34677(.A (u6_mem_b3_b_141 ), .B (n_7758), .Y (n_7747));
NAND2X1 g34676(.A (u6_mem_b3_b_122 ), .B (n_7758), .Y (n_7748));
NAND2X1 g34675(.A (u6_mem_b3_b_140 ), .B (n_7758), .Y (n_7749));
NAND2X1 g34674(.A (u6_mem_b3_b_139 ), .B (n_7758), .Y (n_7750));
OAI21X1 g33953(.A0 (n_4272), .A1 (n_8898), .B0 (n_7574), .Y (n_8875));
NAND2X1 g34672(.A (u6_mem_b3_b_137 ), .B (n_7758), .Y (n_7752));
OAI21X1 g33951(.A0 (n_4497), .A1 (n_8898), .B0 (n_7576), .Y (n_8878));
NAND2X1 g34670(.A (u6_mem_b3_b_135 ), .B (n_7758), .Y (n_7754));
NAND2X1 g34679(.A (u6_mem_b3_b_143 ), .B (n_7758), .Y (n_7745));
NAND2X1 g34678(.A (u6_mem_b3_b_142 ), .B (n_7758), .Y (n_7746));
MX2X1 g38704(.A (u7_mem_b0_b_107 ), .B (wb_din_677), .S0 (n_3622), .Y(n_3644));
AOI22X1 g37923(.A0 (u10_din_tmp_43), .A1 (n_3339), .B0 (n_3911), .B1(in_slt_422), .Y (n_4559));
NAND2X1 g39623(.A (u5_mem_b2_b_44 ), .B (n_12823), .Y (n_11967));
NAND2X1 g39622(.A (u6_mem_b1_b_89 ), .B (n_12169), .Y (n_4159));
NAND2X1 g39621(.A (u6_mem_b2_b_58 ), .B (n_3423), .Y (n_3054));
NAND2X1 g39620(.A (n_4560), .B (in_slt_455), .Y (n_5307));
NAND2X1 g39627(.A (u6_mem_b2_b_59 ), .B (n_3423), .Y (n_3051));
NAND2X1 g39626(.A (u8_mem_b2_b_48 ), .B (n_3441), .Y (n_3052));
NAND2X1 g39625(.A (u6_mem_b2_b_46 ), .B (n_2285), .Y (n_2274));
NAND2X1 g39624(.A (u6_mem_b1_b_77 ), .B (n_4253), .Y (n_4158));
NAND2X1 g39629(.A (u6_mem_b1_b_78 ), .B (n_12169), .Y (n_4157));
MX2X1 g38703(.A (u7_mem_b0_b_105 ), .B (wb_din_675), .S0 (n_3622), .Y(n_3645));
NAND2X1 g34453(.A (u4_mem_b3_b_143 ), .B (n_7984), .Y (n_7968));
OAI21X1 g33480(.A0 (n_5134), .A1 (n_8375), .B0 (n_8091), .Y (n_8376));
NAND2X1 g34451(.A (n_6042), .B (n_7442), .Y (n_7515));
OAI21X1 g33482(.A0 (n_4958), .A1 (n_8372), .B0 (n_8088), .Y (n_8373));
OAI21X1 g33485(.A0 (n_5120), .A1 (n_8372), .B0 (n_8063), .Y (n_8368));
NAND2X1 g34456(.A (u4_mem_b3_b_146 ), .B (n_7984), .Y (n_7965));
NAND2X1 g34455(.A (u4_mem_b3_b_145 ), .B (n_7984), .Y (n_7966));
OR2X1 g34902(.A (n_7434), .B (n_11534), .Y (n_7519));
OAI21X1 g33489(.A0 (n_5142), .A1 (n_8369), .B0 (n_8083), .Y (n_8364));
OAI21X1 g33488(.A0 (n_3887), .A1 (n_8894), .B0 (n_8080), .Y (n_8365));
NAND2X1 g34459(.A (u4_mem_b3_b_149 ), .B (n_7984), .Y (n_7962));
NAND2X1 g34458(.A (u4_mem_b3_b_148 ), .B (n_7984), .Y (n_7963));
MX2X1 g34909(.A (i3_full), .B (u14_u6_full_empty_r), .S0 (n_7389), .Y(n_8215));
NOR2X1 g41405(.A (n_8536), .B (oc3_cfg_997), .Y (n_9656));
NAND2X1 g41407(.A (u13_intm_r_b0_b ), .B (u13_ints_r_b0_b ), .Y(n_442));
NOR2X1 g39842(.A (n_3486), .B (n_2702), .Y (n_2928));
AND2X1 g41401(.A (n_590), .B (n_127), .Y (n_9717));
INVX1 g45563(.A (n_12167), .Y (n_12172));
BUFX3 g41151(.A (n_1147), .Y (n_5112));
NAND2X1 g45886(.A (n_12619), .B (u3_mem_b2_b_40 ), .Y (n_12617));
CLKBUFX1 g45880(.A (n_12607), .Y (n_12608));
NAND4X1 g45882(.A (n_12611), .B (n_12612), .C (n_12613), .D(n_12617), .Y (n_12618));
NAND2X1 g45883(.A (n_3316), .B (u3_mem_b1_b_71 ), .Y (n_12611));
AND2X1 g45889(.A (n_600), .B (u3_rp_b2_b ), .Y (n_12614));
NAND2X2 g45562(.A (n_11587), .B (n_782), .Y (n_12167));
AOI21X1 g30026(.A0 (n_9607), .A1 (n_9768), .B0 (n_10401), .Y(n_10809));
NAND2X1 g34435(.A (u4_mem_b3_b_134 ), .B (n_7984), .Y (n_7980));
XOR2X1 g35504(.A (u26_cnt_b0_b ), .B (n_5624), .Y (n_5615));
AOI21X1 g30025(.A0 (n_9557), .A1 (n_9701), .B0 (n_10090), .Y(n_10409));
XOR2X1 g35502(.A (n_5616), .B (n_4090), .Y (n_5617));
AOI21X1 g35503(.A0 (u11_rp_b0_b ), .A1 (i6_re), .B0 (n_6709), .Y(n_7141));
AND2X1 g30020(.A (n_11151), .B (n_991), .Y (n_11165));
NAND2X1 g34434(.A (u4_mem_b3_b_133 ), .B (n_7984), .Y (n_7981));
AND2X1 g38909(.A (n_869), .B (wb_cyc_i), .Y (n_1284));
NAND2X1 g34437(.A (u4_mem_b3_b_136 ), .B (n_7984), .Y (n_7978));
AOI21X1 g30028(.A0 (n_9605), .A1 (n_9766), .B0 (n_10400), .Y(n_10808));
AOI21X1 g30029(.A0 (n_9553), .A1 (n_9697), .B0 (n_10088), .Y(n_10407));
NAND2X1 g34436(.A (u4_mem_b3_b_135 ), .B (n_7984), .Y (n_7979));
INVX2 g41158(.A (n_1409), .Y (n_2736));
NAND2X1 g34430(.A (u4_mem_b3_b ), .B (n_7984), .Y (n_7986));
OAI21X1 g33688(.A0 (n_4978), .A1 (n_9212), .B0 (n_7851), .Y (n_9211));
OAI21X1 g33425(.A0 (n_3888), .A1 (n_8464), .B0 (n_8153), .Y (n_8443));
NAND2X1 g38908(.A (u3_mem_b3_b_127 ), .B (n_1517), .Y (n_1532));
AOI21X1 g35626(.A0 (n_6300), .A1 (n_6094), .B0 (n_12640), .Y(n_7241));
OAI21X1 g33424(.A0 (n_5150), .A1 (n_8440), .B0 (n_8058), .Y (n_8445));
INVX1 g42171(.A (u11_mem_b3_b_62 ), .Y (n_6658));
NAND2X1 g34349(.A (u4_mem_b1_b_69 ), .B (n_7984), .Y (n_8055));
MX2X1 g38637(.A (u4_mem_b0_b_97 ), .B (wb_din_667), .S0 (n_3765), .Y(n_3754));
NAND2X1 g34348(.A (u4_mem_b1_b ), .B (n_7984), .Y (n_8056));
INVX1 g42172(.A (u10_mem_b3_b_87 ), .Y (n_5504));
MX2X1 g38635(.A (u4_mem_b0_b_94 ), .B (wb_din_664), .S0 (n_3765), .Y(n_3756));
NAND2X1 g34714(.A (u3_mem_b2_b_44 ), .B (n_8141), .Y (n_7723));
MX2X1 g38634(.A (u4_mem_b0_b_93 ), .B (wb_din_663), .S0 (n_3765), .Y(n_3757));
AOI21X1 g38170(.A0 (u4_mem_b2_b_30 ), .A1 (n_4439), .B0 (n_2205), .Y(n_4418));
AOI21X1 g38171(.A0 (u4_mem_b2_b_58 ), .A1 (n_4439), .B0 (n_2478), .Y(n_4417));
AOI21X1 g38172(.A0 (u4_mem_b2_b_59 ), .A1 (n_4439), .B0 (n_1632), .Y(n_4416));
AOI21X1 g38173(.A0 (u6_mem_b2_b_36 ), .A1 (n_4544), .B0 (n_2089), .Y(n_4415));
AOI21X1 g38174(.A0 (u4_mem_b2_b_31 ), .A1 (n_4439), .B0 (n_2206), .Y(n_4414));
NAND2X1 g34864(.A (u3_mem_b1_b_81 ), .B (n_8141), .Y (n_7570));
AOI21X1 g38176(.A0 (u8_mem_b1_b ), .A1 (n_4502), .B0 (n_2091), .Y(n_4412));
AOI21X1 g38177(.A0 (u4_mem_b2_b_33 ), .A1 (n_4439), .B0 (n_2077), .Y(n_4411));
NAND2X1 g34865(.A (u8_mem_b2_b_51 ), .B (n_7976), .Y (n_7569));
MX2X1 g38631(.A (u4_mem_b0_b_92 ), .B (wb_din_662), .S0 (n_835), .Y(n_3761));
NAND2X1 g34710(.A (n_7441), .B (n_7439), .Y (n_8208));
MX2X1 g38630(.A (u4_mem_b0_b_119 ), .B (wb_din_689), .S0 (n_3765), .Y(n_3762));
NAND2X1 g39845(.A (n_12839), .B (u4_mem_b0_b_118 ), .Y (n_2926));
NAND2X1 g34863(.A (u8_mem_b2_b_49 ), .B (n_7976), .Y (n_7571));
NOR2X1 g40137(.A (n_2784), .B (n_2729), .Y (n_2754));
NOR2X1 g40135(.A (n_2099), .B (n_2684), .Y (n_2100));
NOR2X1 g40134(.A (n_2732), .B (n_2137), .Y (n_2176));
NOR2X1 g40133(.A (n_2171), .B (n_2864), .Y (n_2172));
NOR2X1 g40132(.A (n_2477), .B (n_2720), .Y (n_2102));
NOR2X1 g40131(.A (n_2103), .B (n_2790), .Y (n_2104));
NOR2X1 g40130(.A (n_945), .B (n_2801), .Y (n_2105));
NAND2X1 g34713(.A (u3_mem_b2_b_29 ), .B (n_8101), .Y (n_7724));
NOR2X1 g40139(.A (n_1147), .B (n_2744), .Y (n_2753));
NOR2X1 g40138(.A (n_2096), .B (n_2681), .Y (n_2097));
AOI21X1 g38282(.A0 (u4_mem_b1_b_69 ), .A1 (n_4471), .B0 (n_2142), .Y(n_4381));
AOI21X1 g38283(.A0 (u5_mem_b1_b_82 ), .A1 (n_5048), .B0 (n_2685), .Y(n_5029));
AOI21X1 g38280(.A0 (u5_mem_b1_b_80 ), .A1 (n_5037), .B0 (n_2754), .Y(n_5031));
AOI21X1 g38281(.A0 (u5_mem_b1_b_81 ), .A1 (n_5048), .B0 (n_2667), .Y(n_5030));
AOI21X1 g38286(.A0 (u5_mem_b1_b_85 ), .A1 (n_5048), .B0 (n_2665), .Y(n_5026));
AOI21X1 g38287(.A0 (u5_mem_b1_b_86 ), .A1 (n_5037), .B0 (n_2823), .Y(n_5025));
AOI21X1 g38284(.A0 (u5_mem_b1_b_83 ), .A1 (n_5048), .B0 (n_2669), .Y(n_5028));
AOI21X1 g38285(.A0 (u5_mem_b1_b_84 ), .A1 (n_5037), .B0 (n_2771), .Y(n_5027));
AOI21X1 g38288(.A0 (u5_mem_b1_b_87 ), .A1 (n_5037), .B0 (n_2808), .Y(n_5024));
MX2X1 g38639(.A (u4_mem_b0_b_99 ), .B (wb_din_669), .S0 (n_3765), .Y(n_3752));
MX2X1 g38638(.A (u4_mem_b0_b_98 ), .B (wb_din_668), .S0 (n_3765), .Y(n_3753));
MX2X1 g38709(.A (u7_mem_b0_b_116 ), .B (wb_din_686), .S0 (n_3622), .Y(n_3638));
INVX2 g41290(.A (n_604), .Y (n_2502));
NAND2X1 g36578(.A (n_6184), .B (n_12115), .Y (n_6185));
NOR2X1 g41292(.A (u4_rp_b3_b ), .B (u4_wp_b2_b ), .Y (n_441));
MX2X1 g38708(.A (u7_mem_b0_b_114 ), .B (wb_din_684), .S0 (n_3622), .Y(n_3639));
INVX4 g42286(.A (n_6821), .Y (n_784));
AOI22X1 g37346(.A0 (n_4729), .A1 (n_4711), .B0 (n_5591), .B1(n_4710), .Y (n_4712));
AOI22X1 g37347(.A0 (n_5272), .A1 (u13_intm_r_b4_b ), .B0 (n_5277), .B1(crac_din_695), .Y (n_5265));
AOI22X1 g37345(.A0 (n_5272), .A1 (u13_intm_r_b3_b ), .B0 (n_5277), .B1(crac_din_694), .Y (n_5266));
AOI22X1 g37342(.A0 (n_5272), .A1 (u13_intm_r_b2_b ), .B0 (n_5277), .B1(crac_din_693), .Y (n_5270));
AOI22X1 g37343(.A0 (n_4729), .A1 (n_4714), .B0 (n_5591), .B1(n_4713), .Y (n_4715));
AOI22X1 g37340(.A0 (n_5272), .A1 (u13_intm_r_b27_b ), .B0 (n_6972),.B1 (oc3_cfg_996), .Y (n_5273));
AOI22X1 g37341(.A0 (n_5272), .A1 (u13_intm_r_b28_b ), .B0 (n_6972),.B1 (oc3_cfg_997), .Y (n_4716));
AOI22X1 g37838(.A0 (n_6448), .A1 (n_1575), .B0 (n_6524), .B1(n_1831), .Y (n_1587));
AOI22X1 g37839(.A0 (n_1756), .A1 (n_1585), .B0 (n_1584), .B1(n_1643), .Y (n_1586));
AOI22X1 g37348(.A0 (n_4729), .A1 (n_8190), .B0 (n_5591), .B1(n_4708), .Y (n_4709));
AOI22X1 g37349(.A0 (n_5591), .A1 (n_4706), .B0 (n_6972), .B1(oc2_cfg_986), .Y (n_4707));
MX2X1 g33104(.A (n_112), .B (wb_din_669), .S0 (n_8643), .Y (n_8636));
MX2X1 g33105(.A (crac_out_861), .B (wb_din_676), .S0 (n_8643), .Y(n_8635));
MX2X1 g33106(.A (crac_out_863), .B (wb_din_678), .S0 (n_8643), .Y(n_8634));
MX2X1 g33107(.A (crac_out_862), .B (wb_din_677), .S0 (n_8643), .Y(n_8633));
MX2X1 g33100(.A (n_311), .B (wb_din_665), .S0 (n_8643), .Y (n_8640));
MX2X1 g33101(.A (n_149), .B (wb_din_666), .S0 (n_8643), .Y (n_8639));
MX2X1 g33102(.A (n_357), .B (wb_din_667), .S0 (n_8643), .Y (n_8638));
MX2X1 g33103(.A (n_231), .B (wb_din_668), .S0 (n_8643), .Y (n_8637));
NOR2X1 g41558(.A (u5_rp_b3_b ), .B (u5_wp_b2_b ), .Y (n_412));
NOR2X1 g41559(.A (n_742), .B (n_703), .Y (n_1281));
MX2X1 g33108(.A (crac_out_864), .B (wb_din_679), .S0 (n_8643), .Y(n_8631));
MX2X1 g33109(.A (crac_out_865), .B (wb_din_680), .S0 (n_8643), .Y(n_8630));
CLKBUFX3 g45601(.A (n_12273), .Y (n_12261));
NAND2X1 g38900(.A (u6_mem_b3_b_125 ), .B (n_2419), .Y (n_2413));
NAND2X1 g39357(.A (u4_mem_b2_b_40 ), .B (n_12079), .Y (n_3248));
CLKBUFX1 g45606(.A (n_12273), .Y (n_12272));
INVX4 g41103(.A (n_1297), .Y (n_7187));
INVX4 g45607(.A (n_11844), .Y (n_12273));
MX2X1 g31168(.A (n_6580), .B (n_6578), .S0 (n_10565), .Y (n_10567));
MX2X1 g31169(.A (n_6577), .B (n_6575), .S0 (n_10565), .Y (n_10566));
MX2X1 g31164(.A (n_6587), .B (n_6585), .S0 (n_9676), .Y (n_10226));
MX2X1 g31165(.A (n_6015), .B (n_6013), .S0 (n_9676), .Y (n_10225));
MX2X1 g31166(.A (n_6012), .B (n_6010), .S0 (n_10137), .Y (n_10224));
MX2X1 g31167(.A (n_6009), .B (n_6007), .S0 (n_10137), .Y (n_10223));
MX2X1 g31160(.A (n_6600), .B (n_6598), .S0 (n_10137), .Y (n_10232));
MX2X1 g31161(.A (n_6597), .B (n_6595), .S0 (n_10137), .Y (n_10230));
MX2X1 g31162(.A (n_6593), .B (n_6591), .S0 (n_9676), .Y (n_10229));
NAND2X1 g38817(.A (u4_mem_b3_b_122 ), .B (n_4258), .Y (n_4259));
NAND2X1 g38816(.A (u4_mem_b3_b_140 ), .B (n_12744), .Y (n_4260));
OAI21X1 g35889(.A0 (n_5554), .A1 (n_7187), .B0 (n_6789), .Y (n_7193));
OAI21X1 g35888(.A0 (n_5705), .A1 (n_7077), .B0 (n_6236), .Y (n_7095));
INVX1 g42578(.A (u9_mem_b1_b_135 ), .Y (n_6954));
OAI21X1 g35883(.A0 (n_5708), .A1 (n_6995), .B0 (n_5861), .Y (n_7099));
NAND2X1 g38813(.A (u4_mem_b3_b_151 ), .B (n_3556), .Y (n_2607));
OAI21X1 g35881(.A0 (n_5710), .A1 (n_6995), .B0 (n_5871), .Y (n_7100));
OAI21X1 g35880(.A0 (n_5711), .A1 (n_7115), .B0 (n_5873), .Y (n_7101));
OAI21X1 g35887(.A0 (n_5717), .A1 (n_7115), .B0 (n_6240), .Y (n_7116));
OAI21X1 g35886(.A0 (n_5720), .A1 (n_7115), .B0 (n_5858), .Y (n_7096));
OAI21X1 g35885(.A0 (n_5708), .A1 (n_7115), .B0 (n_6143), .Y (n_7047));
AOI21X1 g38192(.A0 (u7_mem_b2_b ), .A1 (n_4540), .B0 (n_2044), .Y(n_4404));
NAND2X1 g38902(.A (u6_mem_b3_b_141 ), .B (n_2465), .Y (n_2411));
NAND2X1 g38811(.A (u4_mem_b3_b_147 ), .B (n_3556), .Y (n_3554));
AOI21X1 g38441(.A0 (u8_mem_b2_b ), .A1 (n_4499), .B0 (n_2092), .Y(n_4328));
NAND2X1 g38810(.A (u4_mem_b3_b_150 ), .B (n_3556), .Y (n_3555));
AOI21X1 g38442(.A0 (u6_mem_b3_b_135 ), .A1 (n_5100), .B0 (n_3333), .Y(n_4924));
AOI21X1 g38196(.A0 (u4_mem_b3_b_138 ), .A1 (n_5102), .B0 (n_3302), .Y(n_5095));
INVX1 g35086(.A (n_7408), .Y (n_9235));
BUFX3 g35084(.A (o4_we), .Y (n_7414));
INVX1 g35088(.A (n_7408), .Y (n_9212));
NOR2X1 g39924(.A (n_3089), .B (n_2804), .Y (n_2873));
INVX1 g42574(.A (u11_mem_b1_b_129 ), .Y (n_6517));
BUFX3 g41560(.A (n_5138), .Y (n_5133));
NAND2X1 g38907(.A (n_685), .B (n_908), .Y (n_4633));
NOR2X1 g39703(.A (n_5102), .B (n_2686), .Y (n_3007));
NOR2X1 g35269(.A (n_7145), .B (n_11597), .Y (n_7372));
NOR2X1 g35268(.A (n_7146), .B (n_11762), .Y (n_7373));
NOR2X1 g35267(.A (n_7147), .B (n_11563), .Y (n_7374));
NOR2X1 g35266(.A (n_7153), .B (n_11762), .Y (n_7375));
NOR2X1 g35265(.A (n_7150), .B (n_11597), .Y (n_7376));
NOR2X1 g35264(.A (n_7152), .B (n_11563), .Y (n_7377));
INVX2 g40730(.A (n_2364), .Y (n_2530));
NAND2X1 g38906(.A (u6_mem_b3_b_139 ), .B (n_2419), .Y (n_2407));
NAND2X1 g39709(.A (n_11789), .B (u8_mem_b0_b_107 ), .Y (n_11668));
INVX1 g42394(.A (oc2_cfg), .Y (n_447));
INVX1 g42397(.A (u10_mem_b0_b_179 ), .Y (n_1251));
INVX2 g42391(.A (n_997), .Y (n_2485));
INVX1 g42390(.A (n_2485), .Y (n_9833));
INVX1 g42392(.A (n_447), .Y (n_997));
NAND2X1 g39164(.A (u7_mem_b1_b_83 ), .B (n_4130), .Y (n_4222));
NAND2X1 g39165(.A (in_slt_407), .B (n_4623), .Y (n_4220));
NAND2X1 g39166(.A (n_11798), .B (u8_mem_b0_b_98 ), .Y (n_11447));
NOR2X1 g39167(.A (n_3453), .B (n_2707), .Y (n_3409));
NAND2X1 g39160(.A (n_6044), .B (n_1300), .Y (n_1453));
NAND2X1 g39161(.A (u3_mem_b1_b_79 ), .B (n_3316), .Y (n_3411));
NOR2X1 g39162(.A (n_2729), .B (n_1488), .Y (n_1492));
NOR2X1 g39163(.A (n_3332), .B (n_2741), .Y (n_3410));
INVX2 g40582(.A (wb_din_661), .Y (n_2707));
INVX1 g43041(.A (n_1873), .Y (n_5827));
NOR2X1 g39168(.A (n_3453), .B (n_2732), .Y (n_3407));
NAND2X1 g39169(.A (n_12826), .B (u3_mem_b0_b_117 ), .Y (n_3406));
INVX1 g43044(.A (oc3_cfg), .Y (n_422));
INVX1 g43045(.A (u9_mem_b0_b_176 ), .Y (n_1728));
INVX2 g32822(.A (n_9737), .Y (n_10277));
NOR2X1 g36829(.A (n_5733), .B (n_5371), .Y (n_5569));
MX2X1 g34028(.A (u5_mem_b0_b_112 ), .B (n_3717), .S0 (n_7496), .Y(n_9424));
MX2X1 g34029(.A (u5_mem_b0_b_113 ), .B (n_3715), .S0 (n_7496), .Y(n_8795));
MX2X1 g34022(.A (u5_mem_b0_b_107 ), .B (n_3728), .S0 (n_7496), .Y(n_8803));
MX2X1 g34023(.A (u5_mem_b0_b_108 ), .B (n_3727), .S0 (n_7496), .Y(n_8801));
MX2X1 g34020(.A (u5_mem_b0_b_105 ), .B (n_3732), .S0 (n_7496), .Y(n_8804));
MX2X1 g34021(.A (u5_mem_b0_b_106 ), .B (n_3731), .S0 (n_7496), .Y(n_9427));
MX2X1 g34026(.A (u5_mem_b0_b_110 ), .B (n_3722), .S0 (n_7496), .Y(n_8798));
MX2X1 g34027(.A (u5_mem_b0_b_111 ), .B (n_3719), .S0 (n_7496), .Y(n_8796));
MX2X1 g34024(.A (u5_mem_b0_b_109 ), .B (n_3725), .S0 (n_7496), .Y(n_9426));
MX2X1 g34025(.A (u5_mem_b0_b_91 ), .B (n_3724), .S0 (n_7496), .Y(n_8800));
AOI21X1 g38092(.A0 (u8_mem_b3_b_142 ), .A1 (n_3879), .B0 (n_1492), .Y(n_3874));
NAND2X1 g36793(.A (n_1767), .B (n_1750), .Y (n_4058));
AOI22X1 g37649(.A0 (n_6931), .A1 (n_1835), .B0 (n_6895), .B1(n_1760), .Y (n_1711));
AOI22X1 g37648(.A0 (n_6888), .A1 (n_1835), .B0 (n_6890), .B1(n_1760), .Y (n_1712));
MX2X1 g38619(.A (u4_mem_b0_b_109 ), .B (wb_din_679), .S0 (n_3765), .Y(n_3783));
NAND2X1 g37138(.A (n_4558), .B (n_1901), .Y (n_6576));
AOI21X1 g38349(.A0 (u6_mem_b3_b_133 ), .A1 (n_5100), .B0 (n_2987), .Y(n_4988));
AOI21X1 g38348(.A0 (u5_mem_b3_b_140 ), .A1 (n_5000), .B0 (n_3132), .Y(n_4989));
AOI21X1 g38347(.A0 (u5_mem_b3_b_139 ), .A1 (n_4996), .B0 (n_2965), .Y(n_4990));
NOR2X1 g37134(.A (n_4268), .B (n_12079), .Y (n_6328));
NAND2X1 g37137(.A (n_4854), .B (n_1411), .Y (n_7049));
NAND2X1 g37136(.A (n_4266), .B (n_12656), .Y (n_6842));
NAND4X1 g37131(.A (n_11449), .B (n_11450), .C (n_2846), .D (n_2370),.Y (n_6260));
INVX1 g37130(.A (n_6260), .Y (n_5667));
NAND2X1 g37133(.A (n_4267), .B (n_2488), .Y (n_6839));
NAND2X1 g37132(.A (n_4269), .B (n_1549), .Y (n_6836));
OAI21X1 g33739(.A0 (n_4476), .A1 (n_9182), .B0 (n_7789), .Y (n_9145));
OAI21X1 g33738(.A0 (n_4468), .A1 (n_9182), .B0 (n_7790), .Y (n_9147));
OAI21X1 g33732(.A0 (n_4934), .A1 (n_9170), .B0 (n_7797), .Y (n_9153));
OAI21X1 g33731(.A0 (n_5108), .A1 (n_9161), .B0 (n_7798), .Y (n_9155));
OAI21X1 g33730(.A0 (n_5097), .A1 (n_9161), .B0 (n_7799), .Y (n_9156));
OAI21X1 g33737(.A0 (n_4338), .A1 (n_9170), .B0 (n_7792), .Y (n_9148));
OAI21X1 g33736(.A0 (n_4443), .A1 (n_9161), .B0 (n_7793), .Y (n_9149));
OAI21X1 g33735(.A0 (n_4906), .A1 (n_9161), .B0 (n_7794), .Y (n_9150));
OAI21X1 g33734(.A0 (n_5111), .A1 (n_9161), .B0 (n_7795), .Y (n_9151));
INVX1 g42408(.A (u9_mem_b0_b_164 ), .Y (n_6396));
INVX1 g42803(.A (u9_mem_b1_b_121 ), .Y (n_6947));
INVX1 g42802(.A (u5_wp_b2_b ), .Y (n_116));
INVX1 g42808(.A (u10_mem_b0_b_168 ), .Y (n_337));
NOR2X1 g40090(.A (n_2775), .B (n_2765), .Y (n_2776));
NOR2X1 g40091(.A (n_945), .B (n_2765), .Y (n_2141));
NOR2X1 g40092(.A (n_2773), .B (n_2772), .Y (n_2774));
NOR2X1 g40093(.A (n_2770), .B (n_2831), .Y (n_2771));
NOR2X1 g40094(.A (n_2470), .B (n_2782), .Y (n_2140));
AOI21X1 g40095(.A0 (oc0_cfg_964), .A1 (in_slt_753), .B0(u14_u0_full_empty_r), .Y (n_635));
NOR2X1 g40096(.A (n_1016), .B (n_2767), .Y (n_2769));
NOR2X1 g40097(.A (n_3008), .B (n_2137), .Y (n_2138));
NOR2X1 g40098(.A (n_2135), .B (n_2829), .Y (n_2136));
NOR2X1 g40099(.A (n_2751), .B (n_2765), .Y (n_2766));
NAND2X1 g36518(.A (n_6816), .B (n_5837), .Y (n_5838));
NAND2X1 g36519(.A (n_6816), .B (n_5835), .Y (n_5836));
INVX4 g40589(.A (wb_din), .Y (n_2801));
NAND2X1 g36510(.A (n_6783), .B (n_6816), .Y (n_6784));
NAND2X1 g36511(.A (n_6228), .B (n_6773), .Y (n_6229));
NAND2X1 g36513(.A (n_6226), .B (n_6816), .Y (n_6227));
NAND2X1 g36514(.A (n_6224), .B (n_1297), .Y (n_6225));
NAND2X1 g36515(.A (n_12368), .B (n_784), .Y (n_6223));
NAND2X1 g36516(.A (n_6816), .B (n_5841), .Y (n_5842));
NOR2X1 g36517(.A (o3_status), .B (n_5839), .Y (n_5840));
INVX1 g42948(.A (u9_mem_b3_b_70 ), .Y (n_6505));
INVX1 g42949(.A (u15_rdd3), .Y (n_294));
INVX1 g42940(.A (u11_mem_b0_b_173 ), .Y (n_1615));
NAND2X1 g45662(.A (n_12531), .B (n_12354), .Y (n_12355));
INVX1 g42945(.A (u11_mem_b2_b_118 ), .Y (n_122));
INVX1 g42947(.A (u9_mem_b1_b_144 ), .Y (n_1703));
INVX1 g40899(.A (n_2553), .Y (n_1232));
INVX4 g40603(.A (wb_din_672), .Y (n_2829));
NAND2X1 g40894(.A (n_403), .B (n_5420), .Y (n_1164));
INVX2 g40897(.A (n_1232), .Y (n_2534));
NAND2X1 g36777(.A (n_1258), .B (wb_addr_i_b6_b), .Y (n_2610));
INVX1 g36770(.A (o8_status), .Y (n_5394));
INVX1 g36773(.A (o9_status), .Y (n_4068));
AND2X1 g41763(.A (n_744), .B (n_444), .Y (n_835));
NAND2X1 g36778(.A (n_1258), .B (n_2608), .Y (n_2609));
AND2X1 g36779(.A (n_1277), .B (u2_res_cnt_b2_b ), .Y (n_1278));
INVX1 g42491(.A (u10_mem_b0_b_169 ), .Y (n_1246));
INVX1 g42494(.A (u10_mem_b2_b_91 ), .Y (n_6630));
INVX1 g42498(.A (u10_mem_b1_b_119 ), .Y (n_406));
NAND3X1 g30912(.A (n_8526), .B (n_8528), .C (n_9498), .Y (n_9525));
NAND3X1 g30913(.A (n_8565), .B (n_8567), .C (n_9559), .Y (n_9601));
AND2X1 g30910(.A (n_9840), .B (n_11564), .Y (n_10335));
NAND3X1 g30916(.A (n_8188), .B (n_8190), .C (n_9496), .Y (n_9523));
NAND3X1 g30917(.A (n_8197), .B (n_8199), .C (n_9495), .Y (n_9522));
NAND3X1 g30914(.A (n_8550), .B (oc2_cfg_987), .C (n_9497), .Y(n_9524));
NAND3X1 g30915(.A (n_8536), .B (oc3_cfg_997), .C (n_9558), .Y(n_9600));
NAND2X1 g39429(.A (n_12389), .B (u4_mem_b0_b_98 ), .Y (n_11660));
NAND2X2 g39428(.A (n_3259), .B (u5_mem_b0_b_95 ), .Y (n_2560));
NOR2X1 g30918(.A (n_9597), .B (u26_ps_cnt_b0_b ), .Y (n_9599));
NOR2X1 g30919(.A (n_1441), .B (n_9597), .Y (n_9598));
INVX1 g41841(.A (wb_addr_i_b4_b), .Y (n_1300));
OAI21X1 g33931(.A0 (n_5144), .A1 (n_8911), .B0 (n_7593), .Y (n_8905));
OAI21X1 g33930(.A0 (n_4393), .A1 (n_8898), .B0 (n_7594), .Y (n_8906));
OAI21X1 g33933(.A0 (n_4402), .A1 (n_8464), .B0 (n_8124), .Y (n_8902));
OAI21X1 g33932(.A0 (n_3841), .A1 (n_8449), .B0 (n_8165), .Y (n_8903));
OAI21X1 g33935(.A0 (n_4503), .A1 (n_8894), .B0 (n_7590), .Y (n_8900));
OAI21X1 g33934(.A0 (n_5143), .A1 (n_8856), .B0 (n_7591), .Y (n_8901));
OAI21X1 g33937(.A0 (n_4913), .A1 (n_8097), .B0 (n_7725), .Y (n_8897));
OAI21X1 g33936(.A0 (n_4302), .A1 (n_8898), .B0 (n_7726), .Y (n_8899));
OAI21X1 g33939(.A0 (n_4275), .A1 (n_8894), .B0 (n_7586), .Y (n_8895));
OAI21X1 g33938(.A0 (n_4274), .A1 (n_8898), .B0 (n_7587), .Y (n_8896));
OAI21X1 g45540(.A0 (n_6078), .A1 (n_11934), .B0 (n_6255), .Y(n_12147));
INVX1 g42239(.A (u10_mem_b1_b_127 ), .Y (n_6037));
MX2X1 g31205(.A (n_6458), .B (n_6457), .S0 (n_10315), .Y (n_10211));
MX2X1 g31204(.A (n_6461), .B (n_6460), .S0 (n_10513), .Y (n_10521));
MX2X1 g31207(.A (n_5979), .B (n_5978), .S0 (n_10839), .Y (n_10841));
MX2X1 g31206(.A (n_5995), .B (n_5994), .S0 (n_10513), .Y (n_10514));
MX2X1 g31201(.A (n_6670), .B (n_461), .S0 (n_10537), .Y (n_10535));
MX2X1 g31200(.A (n_6472), .B (n_6471), .S0 (n_10537), .Y (n_10538));
MX2X1 g31203(.A (n_6464), .B (n_6463), .S0 (n_10315), .Y (n_10212));
MX2X1 g31202(.A (n_6467), .B (n_6466), .S0 (n_10537), .Y (n_10529));
MX2X1 g31209(.A (n_6455), .B (n_6454), .S0 (n_10839), .Y (n_10840));
MX2X1 g31208(.A (n_6536), .B (n_508), .S0 (n_10315), .Y (n_10205));
OAI21X1 g45543(.A0 (n_12156), .A1 (n_12157), .B0 (n_12161), .Y(n_12195));
NAND2X1 g39398(.A (n_12679), .B (u5_mem_b0_b_120 ), .Y (n_3212));
XOR2X1 g40446(.A (n_1203), .B (n_4074), .Y (n_1204));
NAND2X1 g39393(.A (u5_mem_b1_b_88 ), .B (n_3239), .Y (n_3215));
NAND2X1 g39392(.A (u5_mem_b2_b_57 ), .B (n_12823), .Y (n_2312));
NOR2X1 g39390(.A (u9_mem_b2_b ), .B (n_1221), .Y (n_1220));
NAND2X1 g39397(.A (u3_mem_b1_b_80 ), .B (n_3316), .Y (n_3213));
NAND2X1 g39396(.A (n_12261), .B (u4_mem_b1_b_70 ), .Y (n_11476));
NAND2X1 g39395(.A (u5_mem_b2_b_45 ), .B (n_12823), .Y (n_12858));
NAND2X1 g39394(.A (n_12679), .B (u5_mem_b0_b_119 ), .Y (n_3214));
INVX2 g34929(.A (n_7428), .Y (n_9182));
INVX1 g34928(.A (n_7428), .Y (n_9170));
INVX1 g34926(.A (n_7428), .Y (n_9080));
INVX1 g34925(.A (n_7428), .Y (n_9105));
INVX1 g34923(.A (n_7428), .Y (n_9077));
INVX1 g34922(.A (n_7428), .Y (n_9100));
INVX1 g34921(.A (n_7428), .Y (n_9087));
AOI22X1 g35696(.A0 (n_6686), .A1 (i6_dout_628), .B0 (i3_dout_566),.B1 (n_6700), .Y (n_6691));
AOI22X1 g35697(.A0 (n_6686), .A1 (i6_dout_629), .B0 (i3_dout_567),.B1 (n_6700), .Y (n_6688));
AOI22X1 g35694(.A0 (n_6686), .A1 (i6_dout_655), .B0 (i3_dout_593),.B1 (n_6700), .Y (n_6743));
AOI22X1 g35695(.A0 (n_6686), .A1 (i6_dout_656), .B0 (i3_dout_594),.B1 (n_6700), .Y (n_6692));
AOI22X1 g35692(.A0 (n_6686), .A1 (i6_dout_654), .B0 (i3_dout_592),.B1 (n_6700), .Y (n_6737));
AOI22X1 g35693(.A0 (n_6686), .A1 (i6_dout_627), .B0 (i3_dout_565),.B1 (n_6700), .Y (n_6738));
AOI22X1 g35690(.A0 (n_6686), .A1 (i6_dout_652), .B0 (i3_dout_590),.B1 (n_6700), .Y (n_6694));
AOI22X1 g35691(.A0 (n_6686), .A1 (i6_dout_653), .B0 (i3_dout_591),.B1 (n_6700), .Y (n_6693));
CLKBUFX3 g41236(.A (n_839), .Y (n_1517));
AOI22X1 g35698(.A0 (n_6686), .A1 (i6_dout_630), .B0 (i3_dout_568),.B1 (n_6700), .Y (n_6687));
AOI22X1 g35699(.A0 (n_6686), .A1 (i6_dout_631), .B0 (i3_dout_569),.B1 (n_6700), .Y (n_6068));
INVX1 g40762(.A (n_1174), .Y (n_2103));
INVX2 g40763(.A (n_938), .Y (n_1174));
OAI21X1 g33427(.A0 (n_5149), .A1 (n_8440), .B0 (n_8064), .Y (n_8441));
CLKBUFX1 g45861(.A (n_12584), .Y (n_12585));
INVX2 g40561(.A (wb_din_667), .Y (n_2712));
INVX2 g40568(.A (wb_din_666), .Y (n_2765));
INVX1 g40760(.A (n_1174), .Y (n_2020));
NAND2X1 g37184(.A (n_4559), .B (n_2290), .Y (n_6579));
AOI22X1 g37639(.A0 (n_2502), .A1 (n_1728), .B0 (n_1727), .B1(n_1859), .Y (n_1729));
INVX1 g40761(.A (n_1174), .Y (n_2043));
AOI22X1 g37636(.A0 (n_2502), .A1 (n_1733), .B0 (n_1732), .B1(n_1859), .Y (n_1734));
NAND3X1 g37189(.A (n_1553), .B (n_1281), .C (n_4088), .Y (n_2615));
AOI21X1 g38112(.A0 (u6_mem_b2_b_39 ), .A1 (n_4504), .B0 (n_2173), .Y(n_4468));
AOI21X1 g38110(.A0 (u4_mem_b1_b_71 ), .A1 (n_4507), .B0 (n_1792), .Y(n_4470));
AOI21X1 g38111(.A0 (u4_mem_b1_b_72 ), .A1 (n_4507), .B0 (n_2180), .Y(n_4469));
AOI21X1 g38116(.A0 (u4_mem_b1_b_76 ), .A1 (n_4507), .B0 (n_1943), .Y(n_4464));
AOI21X1 g38117(.A0 (u4_mem_b1_b_77 ), .A1 (n_4471), .B0 (n_2151), .Y(n_4463));
AOI21X1 g38115(.A0 (u4_mem_b1_b_74 ), .A1 (n_4507), .B0 (n_1957), .Y(n_4465));
AOI22X1 g37632(.A0 (n_35), .A1 (n_1835), .B0 (n_5374), .B1 (n_1760),.Y (n_1741));
AOI21X1 g38118(.A0 (u4_mem_b1_b_78 ), .A1 (n_4471), .B0 (n_2161), .Y(n_4462));
INVX1 g40766(.A (n_1174), .Y (n_2038));
INVX1 g41741(.A (n_1040), .Y (n_1360));
NAND2X1 g39408(.A (n_3255), .B (u5_mem_b0_b_91 ), .Y (n_3202));
AOI21X1 g30938(.A0 (resume_req), .A1 (suspended_o), .B0(u2_sync_resume), .Y (n_9521));
NOR2X1 g41745(.A (u13_ints_r_b9_b ), .B (n_665), .Y (n_666));
INVX1 g40767(.A (n_1174), .Y (n_2059));
NAND2X1 g41744(.A (n_431), .B (n_667), .Y (n_830));
NOR2X1 g40151(.A (n_2742), .B (n_2741), .Y (n_2743));
NOR2X1 g40150(.A (n_941), .B (n_2772), .Y (n_2089));
NOR2X1 g40153(.A (n_938), .B (n_2691), .Y (n_2087));
NOR2X1 g40152(.A (n_2713), .B (n_2767), .Y (n_2740));
NOR2X1 g40155(.A (n_2083), .B (n_2831), .Y (n_2084));
NOR2X1 g40154(.A (n_2085), .B (n_2864), .Y (n_2086));
NOR2X1 g40157(.A (n_2099), .B (n_2765), .Y (n_2372));
NAND2X1 g39402(.A (u5_mem_b1_b_90 ), .B (n_3209), .Y (n_3210));
NOR2X1 g40159(.A (n_2135), .B (n_2691), .Y (n_2080));
NOR2X1 g40158(.A (n_2784), .B (n_2794), .Y (n_2967));
NAND2X1 g39400(.A (u7_mem_b2_b_44 ), .B (n_12641), .Y (n_4196));
INVX8 g32928(.A (n_9820), .Y (n_10537));
INVX1 g40764(.A (n_1174), .Y (n_2025));
NOR2X1 g39407(.A (n_5059), .B (n_2794), .Y (n_3204));
NOR2X1 g30931(.A (n_9484), .B (n_9587), .Y (n_9588));
NAND2X1 g39405(.A (u5_mem_b1_b_78 ), .B (n_3209), .Y (n_3206));
NAND2X1 g39404(.A (u3_mem_b2_b_38 ), .B (n_3207), .Y (n_3208));
NOR2X1 g39995(.A (n_2171), .B (n_2801), .Y (n_2210));
NOR2X1 g41317(.A (n_4074), .B (u9_wp_b2_b ), .Y (n_1059));
OAI21X1 g33836(.A0 (n_4891), .A1 (n_9055), .B0 (n_7687), .Y (n_9025));
OAI21X1 g33837(.A0 (n_5079), .A1 (n_9034), .B0 (n_7686), .Y (n_9024));
NOR2X1 g37584(.A (n_5321), .B (n_6649), .Y (n_4637));
NOR2X1 g37586(.A (n_5300), .B (n_6649), .Y (n_4635));
OAI21X1 g33918(.A0 (n_4386), .A1 (n_8457), .B0 (n_7604), .Y (n_8924));
NOR2X1 g37580(.A (n_4778), .B (n_5371), .Y (n_3946));
NAND2X1 g37581(.A (n_5645), .B (n_4108), .Y (n_5227));
NAND2X1 g37582(.A (n_3985), .B (n_593), .Y (n_1776));
OAI21X1 g33839(.A0 (n_4890), .A1 (n_9034), .B0 (n_7685), .Y (n_9021));
INVX8 g41313(.A (n_1846), .Y (n_6856));
INVX1 g37588(.A (n_1815), .Y (n_1258));
NOR2X1 g39990(.A (n_2832), .B (n_2831), .Y (n_2833));
OAI21X1 g33694(.A0 (n_4970), .A1 (n_9202), .B0 (n_7845), .Y (n_9204));
OAI21X1 g33695(.A0 (n_4969), .A1 (n_9202), .B0 (n_7844), .Y (n_9203));
OAI21X1 g33696(.A0 (n_4950), .A1 (n_9205), .B0 (n_7843), .Y (n_9201));
OAI21X1 g33697(.A0 (n_4968), .A1 (n_9205), .B0 (n_7842), .Y (n_9200));
OAI21X1 g33690(.A0 (n_4976), .A1 (n_9230), .B0 (n_7849), .Y (n_9209));
OAI21X1 g33691(.A0 (n_4974), .A1 (n_9230), .B0 (n_7848), .Y (n_9208));
OAI21X1 g33692(.A0 (n_4972), .A1 (n_9205), .B0 (n_7847), .Y (n_9207));
OAI21X1 g33693(.A0 (n_4971), .A1 (n_9205), .B0 (n_7846), .Y (n_9206));
OAI21X1 g35941(.A0 (n_5679), .A1 (n_7077), .B0 (n_6168), .Y (n_7059));
OAI21X1 g33698(.A0 (n_4966), .A1 (n_9202), .B0 (n_7841), .Y (n_9199));
AND2X1 g35452(.A (n_4843), .B (u2_sync_resume), .Y (n_5627));
OAI21X1 g33912(.A0 (n_4380), .A1 (n_8930), .B0 (n_7839), .Y (n_8932));
NAND2X1 g38996(.A (u8_mem_b3_b_132 ), .B (n_2468), .Y (n_2373));
OAI21X1 g33911(.A0 (n_4286), .A1 (n_8933), .B0 (n_7611), .Y (n_8934));
OAI21X1 g33910(.A0 (n_4391), .A1 (n_8933), .B0 (n_7612), .Y (n_8935));
NAND2X1 g34637(.A (u6_mem_b2_b_41 ), .B (n_7758), .Y (n_7788));
NAND2X1 g38995(.A (u8_mem_b3_b_142 ), .B (n_2468), .Y (n_2374));
NAND2X1 g38800(.A (u6_mem_b3_b_149 ), .B (n_2465), .Y (n_2458));
AOI22X1 g37361(.A0 (n_5272), .A1 (u13_intm_r_b12_b ), .B0 (n_5277),.B1 (crac_din_703), .Y (n_5255));
AOI22X1 g37362(.A0 (n_5272), .A1 (u13_intm_r_b18_b ), .B0(u13_ints_r_b18_b ), .B1 (n_4726), .Y (n_4694));
AOI22X1 g37363(.A0 (n_4729), .A1 (oc5_cfg_1020), .B0 (n_5591), .B1(ic1_cfg_1040), .Y (n_4693));
AOI22X1 g37364(.A0 (n_5272), .A1 (u13_intm_r_b13_b ), .B0 (n_5277),.B1 (crac_din_704), .Y (n_5254));
NAND2X1 g34635(.A (u6_mem_b2_b_39 ), .B (n_7758), .Y (n_7790));
AOI22X1 g37366(.A0 (n_4729), .A1 (oc5_cfg_1016), .B0 (n_5591), .B1(n_4690), .Y (n_4692));
AOI22X1 g37369(.A0 (n_4729), .A1 (n_4688), .B0 (n_5591), .B1(n_4687), .Y (n_4689));
OAI21X1 g33914(.A0 (n_4383), .A1 (n_8933), .B0 (n_7608), .Y (n_8929));
NOR2X1 g41578(.A (n_568), .B (n_936), .Y (n_569));
NOR2X1 g41574(.A (u13_ints_r_b21_b ), .B (ic0_int_set_719), .Y(n_453));
AOI21X1 g38228(.A0 (u4_mem_b3_b_128 ), .A1 (n_5102), .B0 (n_2810), .Y(n_5067));
NOR2X1 g41576(.A (wb_addr_i_b3_b), .B (wb_addr_i_b4_b), .Y (n_7443));
INVX4 g41571(.A (n_5138), .Y (n_1448));
NOR2X1 g41573(.A (n_627), .B (n_626), .Y (n_743));
XOR2X1 g36189(.A (n_1420), .B (n_1790), .Y (n_4842));
XOR2X1 g36188(.A (n_1425), .B (n_1269), .Y (n_4092));
MX2X1 g36183(.A (n_6335), .B (n_6570), .S0 (n_6341), .Y (n_6336));
MX2X1 g36182(.A (n_6337), .B (n_6573), .S0 (n_6341), .Y (n_6338));
MX2X1 g36181(.A (n_6339), .B (n_6576), .S0 (n_6341), .Y (n_6340));
MX2X1 g36180(.A (n_6342), .B (n_6579), .S0 (n_6341), .Y (n_6343));
XOR2X1 g36187(.A (n_920), .B (n_1294), .Y (n_4093));
MX2X1 g36185(.A (n_6333), .B (n_6563), .S0 (n_6341), .Y (n_6334));
MX2X1 g36184(.A (n_5945), .B (n_6003), .S0 (n_6341), .Y (n_5946));
NAND2X1 g36451(.A (n_5886), .B (n_6141), .Y (n_5887));
NOR2X1 g36450(.A (n_1794), .B (n_1793), .Y (n_4084));
INVX2 g42564(.A (u6_rp_b2_b ), .Y (n_782));
NAND2X1 g36453(.A (n_5882), .B (n_5881), .Y (n_5883));
NAND2X1 g36452(.A (n_5884), .B (n_6141), .Y (n_5885));
NAND2X1 g36455(.A (n_5882), .B (n_5876), .Y (n_5878));
NAND2X1 g36454(.A (n_5879), .B (n_5881), .Y (n_5880));
MX2X1 g36105(.A (n_5978), .B (n_5987), .S0 (n_5312), .Y (n_5979));
MX2X1 g36104(.A (n_6457), .B (n_6592), .S0 (n_6475), .Y (n_6458));
CLKBUFX1 g40807(.A (n_995), .Y (n_5405));
NAND2X1 g38967(.A (u3_mem_b3_b_122 ), .B (n_1517), .Y (n_1512));
NAND2X1 g38913(.A (u8_mem_b3_b_139 ), .B (n_2468), .Y (n_1883));
INVX2 g40802(.A (n_995), .Y (n_1090));
NAND2X1 g38966(.A (u3_mem_b3_b_140 ), .B (n_2463), .Y (n_2392));
INVX8 g35067(.A (n_7984), .Y (n_7499));
INVX8 g40800(.A (n_1090), .Y (n_6502));
NAND2X1 g37989(.A (n_2841), .B (n_2997), .Y (n_5161));
NAND2X1 g38965(.A (u8_mem_b3_b_128 ), .B (n_2468), .Y (n_2393));
INVX1 g42009(.A (u10_mem_b0_b_165 ), .Y (n_5957));
INVX1 g42008(.A (u11_mem_b0_b_165 ), .Y (n_5953));
INVX1 g42007(.A (u9_mem_b0_b ), .Y (n_6868));
INVX1 g42001(.A (dma_req_o_b0_b), .Y (n_271));
INVX1 g42002(.A (u9_mem_b0_b_169 ), .Y (n_1742));
NOR2X1 g39986(.A (n_2218), .B (n_2790), .Y (n_2219));
AOI21X1 g39987(.A0 (oc2_cfg_984), .A1 (in_slt_750), .B0(u14_u2_full_empty_r), .Y (n_531));
NOR2X1 g39984(.A (n_2216), .B (n_2864), .Y (n_2222));
NOR2X1 g39985(.A (n_867), .B (n_2829), .Y (n_2221));
NOR2X1 g39983(.A (n_2827), .B (n_2712), .Y (n_2835));
NOR2X1 g39980(.A (n_2832), .B (n_2786), .Y (n_2839));
NOR2X1 g39981(.A (n_2736), .B (n_2829), .Y (n_2838));
NOR2X1 g39988(.A (n_2216), .B (n_3008), .Y (n_2217));
NOR2X1 g39989(.A (n_2786), .B (n_2067), .Y (n_2215));
NAND2X1 g37452(.A (u13_ints_r_b24_b ), .B (n_4726), .Y (n_2586));
NAND2X1 g37453(.A (u13_ints_r_b26_b ), .B (n_4726), .Y (n_2585));
INVX1 g35202(.A (n_7396), .Y (n_8868));
NAND2X1 g37450(.A (u13_ints_r_b13_b ), .B (n_3979), .Y (n_3978));
INVX1 g35206(.A (n_7396), .Y (n_8898));
NAND2X1 g37451(.A (n_5272), .B (u13_intm_r_b23_b ), .Y (n_3976));
AOI22X1 g37984(.A0 (n_2558), .A1 (n_1864), .B0 (n_1863), .B1(n_2544), .Y (n_1865));
NAND2X1 g38963(.A (u8_mem_b3_b ), .B (n_2468), .Y (n_2395));
NAND2X1 g37457(.A (u13_ints_r_b3_b ), .B (n_3979), .Y (n_3974));
NAND2X1 g37454(.A (u13_ints_r_b27_b ), .B (n_4726), .Y (n_2584));
AOI22X1 g37987(.A0 (n_6471), .A1 (n_1575), .B0 (n_6604), .B1(n_1831), .Y (n_1891));
NAND2X1 g39188(.A (u7_mem_b1_b_80 ), .B (n_11856), .Y (n_4217));
NAND2X1 g39189(.A (u4_mem_b2_b_47 ), .B (n_12079), .Y (n_2348));
NAND2X1 g39186(.A (u4_mem_b2_b_59 ), .B (n_12087), .Y (n_3394));
NAND2X1 g39187(.A (n_12389), .B (u4_mem_b0_b_109 ), .Y (n_3393));
NAND2X1 g39184(.A (u3_mem_b1_b_74 ), .B (n_3316), .Y (n_12833));
NAND2X1 g39185(.A (u3_mem_b2_b_41 ), .B (n_12619), .Y (n_3396));
NAND2X1 g39182(.A (u4_mem_b2_b_56 ), .B (n_12091), .Y (n_3399));
NAND2X1 g39183(.A (n_11804), .B (u8_mem_b0_b_112 ), .Y (n_3398));
NAND2X1 g39181(.A (u4_mem_b2_b_46 ), .B (n_12079), .Y (n_2260));
INVX1 g41161(.A (n_1409), .Y (n_2761));
INVX1 g41905(.A (n_746), .Y (n_411));
NAND2X1 g38803(.A (u3_mem_b3_b_150 ), .B (n_2463), .Y (n_1811));
AOI22X1 g37643(.A0 (n_206), .A1 (n_1859), .B0 (n_5345), .B1 (n_1760),.Y (n_1720));
NAND2X1 g38961(.A (u4_mem_b3_b ), .B (n_12744), .Y (n_4250));
NAND2X1 g38842(.A (u5_mem_b3_b_127 ), .B (n_1543), .Y (n_1327));
INVX1 g41907(.A (n_746), .Y (n_1421));
MX2X1 g34004(.A (u4_mem_b0_b_120 ), .B (n_3760), .S0 (n_7499), .Y(n_8816));
MX2X1 g34005(.A (u4_mem_b0_b_121 ), .B (n_3759), .S0 (n_7499), .Y(n_9434));
MX2X1 g34006(.A (u4_mem_b0_b_93 ), .B (n_3757), .S0 (n_7499), .Y(n_8815));
MX2X1 g34007(.A (u4_mem_b0_b_94 ), .B (n_3756), .S0 (n_7499), .Y(n_9433));
MX2X1 g34001(.A (u4_mem_b0_b_118 ), .B (n_3763), .S0 (n_7499), .Y(n_8820));
MX2X1 g34002(.A (u4_mem_b0_b_119 ), .B (n_3762), .S0 (n_7499), .Y(n_8818));
MX2X1 g34008(.A (u4_mem_b0_b_95 ), .B (n_3790), .S0 (n_7499), .Y(n_8813));
NAND2X1 g34558(.A (u5_mem_b3_b_133 ), .B (n_7870), .Y (n_7868));
NAND2X1 g34559(.A (u5_mem_b3_b_134 ), .B (n_7870), .Y (n_7867));
INVX1 g43064(.A (n_706), .Y (n_473));
INVX1 g43066(.A (n_706), .Y (n_1417));
INVX1 g43060(.A (u10_mem_b3_b_76 ), .Y (n_5520));
INVX1 g43061(.A (u9_mem_b0_b_159 ), .Y (n_6404));
INVX1 g43068(.A (u9_mem_b3_b_86 ), .Y (n_5365));
INVX1 g43069(.A (u11_mem_b3_b_80 ), .Y (n_5496));
NOR2X1 g41318(.A (n_605), .B (n_689), .Y (n_606));
NAND2X1 g38807(.A (u8_mem_b3_b_129 ), .B (n_2468), .Y (n_2455));
AOI21X1 g38388(.A0 (u7_mem_b3_b_128 ), .A1 (n_5145), .B0 (n_3454), .Y(n_4956));
AOI21X1 g38343(.A0 (u5_mem_b3_b_136 ), .A1 (n_5000), .B0 (n_2939), .Y(n_4994));
AOI21X1 g38329(.A0 (u5_mem_b2_b_31 ), .A1 (n_4378), .B0 (n_2152), .Y(n_4355));
AOI21X1 g38328(.A0 (u6_mem_b3_b_149 ), .A1 (n_5100), .B0 (n_3234), .Y(n_5006));
AOI21X1 g38321(.A0 (u5_mem_b2_b_53 ), .A1 (n_4378), .B0 (n_1939), .Y(n_4362));
AOI21X1 g38320(.A0 (u5_mem_b2_b_52 ), .A1 (n_4378), .B0 (n_2049), .Y(n_4363));
AOI21X1 g38323(.A0 (u5_mem_b2_b_55 ), .A1 (n_4370), .B0 (n_1949), .Y(n_4360));
AOI21X1 g38322(.A0 (u5_mem_b2_b_54 ), .A1 (n_4378), .B0 (n_2011), .Y(n_4361));
AOI21X1 g38324(.A0 (u5_mem_b2_b_56 ), .A1 (n_4378), .B0 (n_1951), .Y(n_4359));
AOI21X1 g38327(.A0 (u5_mem_b2_b_59 ), .A1 (n_4370), .B0 (n_2225), .Y(n_4356));
AOI21X1 g38326(.A0 (u5_mem_b2_b_57 ), .A1 (n_4370), .B0 (n_2126), .Y(n_4357));
INVX1 g41939(.A (n_12585), .Y (n_8182));
INVX8 g32891(.A (n_9827), .Y (n_10450));
INVX2 g32898(.A (n_10065), .Y (n_9827));
INVX1 g41863(.A (u10_mem_b2_b_93 ), .Y (n_6612));
NAND2X1 g38791(.A (u6_mem_b3_b_144 ), .B (n_2465), .Y (n_2466));
INVX1 g42827(.A (u11_mem_b3_b_81 ), .Y (n_5492));
INVX1 g42826(.A (u10_mem_b2_b_97 ), .Y (n_6610));
INVX1 g42824(.A (u11_mem_b2_b_109 ), .Y (n_279));
INVX1 g41861(.A (u11_mem_b2_b_92 ), .Y (n_6437));
INVX1 g42822(.A (u8_wp_b2_b ), .Y (n_1446));
INVX1 g37117(.A (n_5800), .Y (n_5529));
NAND4X1 g37116(.A (n_12843), .B (n_11501), .C (n_12844), .D (n_2384),.Y (n_6159));
INVX1 g37115(.A (n_6159), .Y (n_5669));
NAND4X1 g37114(.A (n_11741), .B (n_11499), .C (n_11742), .D (n_2435),.Y (n_6250));
INVX1 g37113(.A (n_6250), .Y (n_5670));
MX2X1 g38632(.A (u4_mem_b0_b_120 ), .B (wb_din_690), .S0 (n_3765), .Y(n_3760));
INVX1 g37111(.A (n_12481), .Y (n_5671));
NAND4X1 g37110(.A (n_2352), .B (n_3890), .C (n_2850), .D (n_1883), .Y(n_6153));
NAND2X1 g37686(.A (n_3552), .B (n_3394), .Y (n_4608));
INVX1 g37119(.A (n_5893), .Y (n_5528));
NAND4X1 g37118(.A (n_11463), .B (n_11464), .C (n_1927), .D (n_2382),.Y (n_5800));
NAND2X1 g36573(.A (n_6144), .B (n_12115), .Y (n_6188));
NAND2X1 g36570(.A (n_12618), .B (n_12115), .Y (n_6193));
NAND2X1 g36571(.A (n_12755), .B (n_12115), .Y (n_6191));
NAND2X1 g36576(.A (n_5813), .B (n_6259), .Y (n_5814));
NAND2X1 g36577(.A (n_5811), .B (n_6259), .Y (n_5812));
NAND2X1 g36574(.A (n_5815), .B (n_6259), .Y (n_5816));
NAND2X1 g36575(.A (n_6186), .B (n_12115), .Y (n_6187));
NAND2X1 g41291(.A (n_53), .B (n_121), .Y (n_604));
NAND2X1 g36579(.A (n_6182), .B (n_6259), .Y (n_6183));
INVX1 g42922(.A (u10_mem_b2_b_103 ), .Y (n_6033));
INVX1 g45603(.A (n_12269), .Y (n_12267));
INVX1 g42920(.A (ic2_cfg_1045), .Y (n_431));
INVX1 g42921(.A (u10_mem_b3_b_60 ), .Y (n_6572));
INVX1 g42925(.A (u9_mem_b0_b_167 ), .Y (n_349));
NAND2X1 g36798(.A (n_1681), .B (n_1741), .Y (n_4054));
NAND2X1 g36799(.A (n_1739), .B (n_1736), .Y (n_4053));
NAND2X1 g36796(.A (n_1747), .B (n_1746), .Y (n_4056));
NAND2X1 g36797(.A (n_1745), .B (n_1743), .Y (n_4055));
NAND2X1 g36794(.A (n_1749), .B (n_1834), .Y (n_4057));
OR2X1 g36795(.A (n_1815), .B (wb_addr_i_b6_b), .Y (n_4837));
NAND2X1 g36792(.A (n_1752), .B (n_1751), .Y (n_4059));
NAND2X1 g37854(.A (n_4165), .B (n_3086), .Y (n_12048));
NAND2X1 g36790(.A (n_1759), .B (n_1758), .Y (n_4061));
NAND2X1 g36791(.A (n_1836), .B (n_1753), .Y (n_4060));
OAI21X1 g33815(.A0 (n_4900), .A1 (n_9055), .B0 (n_7712), .Y (n_9054));
NAND2X1 g39553(.A (n_2325), .B (in_slt_454), .Y (n_2288));
INVX2 g41312(.A (n_1059), .Y (n_1846));
NAND2X1 g36585(.A (n_3563), .B (n_2624), .Y (n_4830));
NOR2X1 g40213(.A (n_2751), .B (n_3008), .Y (n_2715));
INVX1 g41743(.A (n_830), .Y (n_831));
INVX1 g41742(.A (n_830), .Y (n_1040));
NAND2X1 g39409(.A (u5_mem_b2_b_29 ), .B (n_12823), .Y (n_11441));
INVX2 g33316(.A (n_12608), .Y (n_9931));
NAND4X1 g33311(.A (n_6049), .B (n_2646), .C (n_7499), .D (n_1001), .Y(n_9452));
AOI21X1 g30939(.A0 (n_11889), .A1 (n_754), .B0 (n_9962), .Y(n_10773));
BUFX3 g41033(.A (n_821), .Y (n_4471));
BUFX3 g41032(.A (n_821), .Y (n_4507));
AOI21X1 g30934(.A0 (n_12339), .A1 (n_763), .B0 (n_9965), .Y(n_10775));
NAND3X1 g30935(.A (n_12077), .B (n_12256), .C (n_10329), .Y(n_10332));
NAND3X1 g30936(.A (n_12214), .B (n_1908), .C (n_10327), .Y (n_10331));
AOI21X1 g30937(.A0 (n_11891), .A1 (n_762), .B0 (n_9963), .Y(n_10774));
NOR2X1 g30930(.A (n_9547), .B (n_9645), .Y (n_9646));
NOR2X1 g30932(.A (n_9482), .B (n_9585), .Y (n_9586));
AOI21X1 g30933(.A0 (n_11893), .A1 (n_12278), .B0 (n_9966), .Y(n_10776));
INVX1 g42210(.A (u9_mem_b1_b_142 ), .Y (n_1732));
OAI21X1 g33919(.A0 (n_4282), .A1 (n_8457), .B0 (n_7603), .Y (n_8922));
NAND2X1 g34638(.A (u6_mem_b2_b_42 ), .B (n_7758), .Y (n_7787));
INVX1 g42215(.A (u10_mem_b1_b_148 ), .Y (n_196));
INVX1 g42217(.A (u10_mem_b3_b_74 ), .Y (n_5577));
OAI21X1 g33913(.A0 (n_4285), .A1 (n_8930), .B0 (n_7610), .Y (n_8931));
NAND2X1 g34632(.A (u6_mem_b2_b ), .B (n_7758), .Y (n_7793));
NAND2X1 g34631(.A (u6_mem_b1_b_68 ), .B (n_7758), .Y (n_7794));
NAND2X1 g34630(.A (u6_mem_b1_b_67 ), .B (n_7758), .Y (n_7795));
OAI21X1 g33917(.A0 (n_4283), .A1 (n_8891), .B0 (n_7605), .Y (n_8925));
OAI21X1 g33916(.A0 (n_4385), .A1 (n_8868), .B0 (n_7945), .Y (n_8926));
OAI21X1 g33915(.A0 (n_4284), .A1 (n_8933), .B0 (n_7606), .Y (n_8928));
NAND2X1 g34634(.A (u3_mem_b1_b_76 ), .B (n_8101), .Y (n_7791));
INVX1 g42665(.A (u11_mem_b3_b_58 ), .Y (n_6524));
MX2X1 g31229(.A (n_6024), .B (n_6023), .S0 (n_10839), .Y (n_10836));
MX2X1 g31228(.A (n_6420), .B (n_6419), .S0 (n_10537), .Y (n_10456));
MX2X1 g31227(.A (n_6422), .B (n_6421), .S0 (n_10537), .Y (n_10457));
MX2X1 g31226(.A (n_6425), .B (n_6424), .S0 (n_10537), .Y (n_10458));
MX2X1 g31225(.A (n_6605), .B (n_6604), .S0 (n_10537), .Y (n_10459));
MX2X1 g31224(.A (n_6427), .B (n_6426), .S0 (n_10537), .Y (n_10462));
MX2X1 g31223(.A (n_6429), .B (n_6428), .S0 (n_10537), .Y (n_10466));
MX2X1 g31222(.A (n_6555), .B (n_6554), .S0 (n_10537), .Y (n_10472));
MX2X1 g31221(.A (n_5970), .B (n_5969), .S0 (n_10537), .Y (n_10476));
MX2X1 g31220(.A (n_6432), .B (n_6431), .S0 (n_10839), .Y (n_10837));
NAND2X1 g34545(.A (u5_mem_b2_b_30 ), .B (n_7870), .Y (n_7882));
NAND2X1 g34544(.A (u5_mem_b2_b_57 ), .B (n_7870), .Y (n_7883));
INVX1 g45418(.A (ic2_cfg), .Y (n_11777));
MX2X1 g34011(.A (u4_mem_b0_b_98 ), .B (n_3753), .S0 (n_7499), .Y(n_8811));
MX2X1 g34010(.A (u4_mem_b0_b_97 ), .B (n_3754), .S0 (n_7499), .Y(n_9432));
NAND2X1 g34541(.A (u5_mem_b2_b_54 ), .B (n_7870), .Y (n_7886));
NAND2X1 g34540(.A (u5_mem_b2_b_53 ), .B (n_7870), .Y (n_7887));
NOR2X1 g32614(.A (n_8479), .B (n_10940), .Y (n_9468));
INVX8 g34941(.A (o7_we), .Y (n_7758));
INVX1 g45413(.A (n_11762), .Y (n_11772));
NAND2X1 g34542(.A (u5_mem_b2_b_55 ), .B (n_7870), .Y (n_7885));
INVX1 g40661(.A (u2_bit_clk_r), .Y (n_719));
INVX1 g42081(.A (u11_mem_b3_b_70 ), .Y (n_6421));
AOI21X1 g34905(.A0 (n_4844), .A1 (n_2302), .B0 (n_4035), .Y (n_6055));
MX2X1 g38707(.A (u7_mem_b0_b_112 ), .B (wb_din_682), .S0 (n_3622), .Y(n_3641));
INVX8 g35171(.A (n_7651), .Y (n_7493));
MX2X1 g38706(.A (u7_mem_b0_b_110 ), .B (wb_din_680), .S0 (n_913), .Y(n_3642));
MX2X1 g38705(.A (u7_mem_b0_b_109 ), .B (wb_din_679), .S0 (n_3622), .Y(n_2635));
NAND4X1 g37063(.A (n_11719), .B (n_11720), .C (n_3208), .D (n_1513),.Y (n_6235));
NOR2X1 g39982(.A (n_2836), .B (n_2748), .Y (n_2837));
INVX1 g37062(.A (n_6235), .Y (n_5685));
INVX4 g40508(.A (wb_din_684), .Y (n_2790));
AOI22X1 g38781(.A0 (n_12291), .A1 (n_6152), .B0 (n_2567), .B1(n_12278), .Y (n_4269));
MX2X1 g38727(.A (u6_mem_b0_b_114 ), .B (wb_din_684), .S0 (n_3632), .Y(n_3614));
INVX1 g42501(.A (u10_mem_b1_b_131 ), .Y (n_6457));
NOR2X1 g30068(.A (n_1870), .B (n_11518), .Y (n_11175));
NOR2X1 g30069(.A (n_11144), .B (n_11516), .Y (n_11174));
NOR2X1 g30062(.A (n_11043), .B (n_11505), .Y (n_11176));
AND2X1 g30063(.A (n_10971), .B (n_991), .Y (n_11157));
OAI21X1 g30060(.A0 (n_9500), .A1 (n_9585), .B0 (n_9753), .Y(n_10087));
INVX2 g40501(.A (wb_din_678), .Y (n_2720));
AND2X1 g30066(.A (n_9757), .B (n_11119), .Y (n_10083));
AND2X1 g30067(.A (n_10970), .B (n_9833), .Y (n_11155));
AND2X1 g30064(.A (n_9693), .B (n_11119), .Y (n_9846));
AND2X1 g30065(.A (n_9692), .B (n_11119), .Y (n_9845));
NAND2X1 g34497(.A (u5_mem_b1_b_75 ), .B (n_7870), .Y (n_7934));
NAND2X1 g34496(.A (u5_mem_b1_b_74 ), .B (n_7870), .Y (n_7935));
NAND2X1 g34495(.A (u5_mem_b1_b_73 ), .B (n_7870), .Y (n_7936));
NAND2X1 g34494(.A (u5_mem_b1_b_72 ), .B (n_7870), .Y (n_7938));
NAND2X1 g34493(.A (u5_mem_b1_b_71 ), .B (n_7870), .Y (n_7939));
NAND2X1 g34492(.A (u5_mem_b1_b_70 ), .B (n_7870), .Y (n_7941));
NAND2X1 g34491(.A (u5_mem_b1_b_69 ), .B (n_7870), .Y (n_7942));
NAND2X2 g34490(.A (n_1225), .B (n_7442), .Y (n_8202));
NAND4X1 g36891(.A (n_2322), .B (n_3258), .C (n_3256), .D (n_1548), .Y(n_6142));
INVX1 g36890(.A (n_6142), .Y (n_5717));
NAND2X1 g36893(.A (n_1669), .B (n_1711), .Y (n_4033));
NAND2X1 g36892(.A (n_2628), .B (n_1241), .Y (n_4817));
NAND4X1 g36895(.A (n_2337), .B (n_3254), .C (n_3194), .D (n_1326), .Y(n_6239));
INVX1 g36894(.A (n_6239), .Y (n_5716));
NAND2X1 g34499(.A (u5_mem_b1_b_77 ), .B (n_7870), .Y (n_7932));
INVX2 g45593(.A (n_12258), .Y (n_12250));
INVX4 g32791(.A (n_9633), .Y (n_10073));
INVX1 g45596(.A (n_12250), .Y (n_12256));
INVX4 g32794(.A (n_9741), .Y (n_10019));
INVX1 g45598(.A (n_12258), .Y (n_12259));
INVX4 g32799(.A (n_9741), .Y (n_10054));
MX2X1 g31106(.A (n_6653), .B (n_6652), .S0 (n_10315), .Y (n_10301));
INVX1 g35545(.A (i6_full), .Y (n_630));
INVX1 g36899(.A (n_6264), .Y (n_5715));
AOI21X1 g38138(.A0 (u4_mem_b1_b_63 ), .A1 (n_4471), .B0 (n_2109), .Y(n_4447));
AOI21X1 g38139(.A0 (u4_mem_b1_b_64 ), .A1 (n_4471), .B0 (n_2047), .Y(n_4446));
NAND4X1 g36898(.A (n_12853), .B (n_12854), .C (n_12796), .D (n_1325),.Y (n_5882));
AOI21X1 g38134(.A0 (u8_mem_b3_b_140 ), .A1 (n_3879), .B0 (n_1483), .Y(n_3867));
AOI21X1 g38135(.A0 (u4_mem_b1_b_89 ), .A1 (n_4507), .B0 (n_2471), .Y(n_4450));
AOI21X1 g38136(.A0 (u4_mem_b1_b_90 ), .A1 (n_4471), .B0 (n_2123), .Y(n_4449));
AOI21X1 g38137(.A0 (u4_mem_b1_b_62 ), .A1 (n_4471), .B0 (n_2483), .Y(n_4448));
AOI21X1 g38130(.A0 (u4_mem_b1_b_86 ), .A1 (n_4507), .B0 (n_2074), .Y(n_4453));
AOI21X1 g38131(.A0 (u7_mem_b2_b_44 ), .A1 (n_4509), .B0 (n_2168), .Y(n_4452));
AOI21X1 g38132(.A0 (u3_mem_b3_b_124 ), .A1 (n_5138), .B0 (n_2873), .Y(n_5115));
AOI21X1 g38133(.A0 (u4_mem_b1_b_61 ), .A1 (n_4507), .B0 (n_2140), .Y(n_4451));
OAI21X1 g36629(.A0 (n_12849), .A1 (n_12850), .B0 (u4_rp_b0_b ), .Y(n_6130));
NOR2X1 g40178(.A (n_2681), .B (n_1985), .Y (n_2292));
NOR2X1 g40173(.A (n_2470), .B (n_2729), .Y (n_2063));
NOR2X1 g40172(.A (n_2020), .B (n_2716), .Y (n_2064));
NOR2X1 g40171(.A (n_2470), .B (n_2786), .Y (n_2065));
NOR2X1 g40170(.A (n_2477), .B (n_2794), .Y (n_2066));
NOR2X1 g40177(.A (n_2736), .B (n_2735), .Y (n_2737));
NOR2X1 g40176(.A (n_2705), .B (n_2794), .Y (n_2738));
NOR2X1 g40175(.A (n_2470), .B (n_2792), .Y (n_2061));
NOR2X1 g40174(.A (n_2684), .B (n_1985), .Y (n_2062));
INVX1 g43078(.A (n_1033), .Y (n_641));
NAND4X1 g36897(.A (n_12032), .B (n_3251), .C (n_12033), .D (n_1542),.Y (n_5884));
NAND2X1 g34498(.A (u5_mem_b1_b_76 ), .B (n_7870), .Y (n_7933));
NAND2X1 g38969(.A (u8_mem_b3_b_133 ), .B (n_2468), .Y (n_2391));
NAND2X1 g38968(.A (u3_mem_b3_b_124 ), .B (n_1517), .Y (n_1511));
NAND2X1 g38790(.A (u3_mem_b3_b_134 ), .B (n_2463), .Y (n_2467));
NAND2X1 g38792(.A (u3_mem_b3_b_151 ), .B (n_2463), .Y (n_2464));
NAND2X1 g38793(.A (u6_mem_b3_b_151 ), .B (n_2465), .Y (n_2462));
NAND2X1 g38794(.A (u3_mem_b3_b_146 ), .B (n_2463), .Y (n_2461));
NAND2X1 g38795(.A (u8_mem_b3_b_144 ), .B (n_2468), .Y (n_2460));
NAND2X1 g37568(.A (n_5645), .B (n_2886), .Y (n_4641));
NOR2X1 g37569(.A (n_4753), .B (n_5371), .Y (n_3948));
NAND2X1 g37566(.A (n_5645), .B (n_4230), .Y (n_5231));
NAND2X1 g37567(.A (n_5645), .B (n_4135), .Y (n_5230));
NAND2X1 g37564(.A (n_5656), .B (n_4209), .Y (n_5233));
NAND2X1 g37565(.A (n_5645), .B (n_4231), .Y (n_5232));
NAND2X1 g37563(.A (n_5656), .B (n_4133), .Y (n_5234));
NAND2X1 g37560(.A (n_5656), .B (n_4207), .Y (n_5237));
NAND2X1 g37561(.A (n_5656), .B (n_4106), .Y (n_5236));
NAND2X1 g38945(.A (u4_mem_b3_b_139 ), .B (n_12744), .Y (n_4252));
INVX1 g42409(.A (u9_mem_b3_b_69 ), .Y (n_6450));
AOI22X1 g37716(.A0 (n_2558), .A1 (n_2557), .B0 (n_2556), .B1(n_2534), .Y (n_2559));
OAI21X1 g33678(.A0 (n_4989), .A1 (n_9205), .B0 (n_7861), .Y (n_9224));
OAI21X1 g33679(.A0 (n_4987), .A1 (n_9205), .B0 (n_7860), .Y (n_9223));
OAI21X1 g33676(.A0 (n_4992), .A1 (n_9205), .B0 (n_7863), .Y (n_9227));
OAI21X1 g33677(.A0 (n_4990), .A1 (n_9205), .B0 (n_7862), .Y (n_9226));
OAI21X1 g33674(.A0 (n_4994), .A1 (n_9230), .B0 (n_7865), .Y (n_9229));
OAI21X1 g33675(.A0 (n_4993), .A1 (n_9230), .B0 (n_7864), .Y (n_9228));
OAI21X1 g33672(.A0 (n_4997), .A1 (n_9230), .B0 (n_7867), .Y (n_9232));
OAI21X1 g33673(.A0 (n_4995), .A1 (n_9230), .B0 (n_7866), .Y (n_9231));
OAI21X1 g33670(.A0 (n_4999), .A1 (n_9235), .B0 (n_7869), .Y (n_9234));
OAI21X1 g33671(.A0 (n_4998), .A1 (n_9235), .B0 (n_7868), .Y (n_9233));
MX2X1 g31810(.A (n_5420), .B (n_5421), .S0 (n_9620), .Y (n_9961));
OAI21X1 g31811(.A0 (n_5634), .A1 (n_9631), .B0 (n_9834), .Y(n_10337));
OAI21X1 g31812(.A0 (n_6056), .A1 (n_9514), .B0 (n_9686), .Y (n_9840));
OAI21X1 g31813(.A0 (n_6055), .A1 (n_9564), .B0 (n_9751), .Y (n_9960));
MX2X1 g31814(.A (u14_u0_full_empty_r), .B (n_9543), .S0 (n_11827), .Y(n_9544));
MX2X1 g31815(.A (u14_u1_full_empty_r), .B (n_9541), .S0 (n_11827), .Y(n_9542));
MX2X1 g31816(.A (u14_u2_full_empty_r), .B (n_9538), .S0 (n_11827), .Y(n_9539));
MX2X1 g31817(.A (u14_u3_full_empty_r), .B (n_9536), .S0 (n_11827), .Y(n_9537));
MX2X1 g31818(.A (u14_u4_full_empty_r), .B (n_9534), .S0 (n_11827), .Y(n_9535));
MX2X1 g31819(.A (u14_u5_full_empty_r), .B (n_9532), .S0 (n_11827), .Y(n_9533));
NAND2X1 g38960(.A (u3_mem_b3_b_147 ), .B (n_2463), .Y (n_2396));
INVX4 g45599(.A (n_12273), .Y (n_12258));
NOR2X1 g39810(.A (n_3089), .B (n_2790), .Y (n_2947));
MX2X1 g37308(.A (u10_mem_b1_b_140 ), .B (n_5290), .S0 (n_6475), .Y(n_5291));
MX2X1 g37309(.A (u10_mem_b1_b_141 ), .B (n_5282), .S0 (n_5407), .Y(n_5289));
NOR2X1 g39811(.A (n_5059), .B (n_2681), .Y (n_2946));
MX2X1 g37302(.A (u11_mem_b2_b_118 ), .B (n_5300), .S0 (n_5409), .Y(n_5301));
MX2X1 g37303(.A (u11_mem_b2_b_116 ), .B (n_5298), .S0 (n_5312), .Y(n_5299));
MX2X1 g37300(.A (u11_mem_b2_b_115 ), .B (n_5304), .S0 (n_5312), .Y(n_5305));
MX2X1 g37306(.A (u10_mem_b1_b_138 ), .B (n_5292), .S0 (n_6475), .Y(n_5293));
MX2X1 g37307(.A (u10_mem_b1_b_139 ), .B (n_4745), .S0 (n_6475), .Y(n_4746));
MX2X1 g37304(.A (u11_mem_b2_b_117 ), .B (n_5296), .S0 (n_5409), .Y(n_5297));
AOI21X1 g37305(.A0 (n_5294), .A1 (n_5371), .B0 (n_3946), .Y (n_5295));
NOR2X1 g39813(.A (n_2686), .B (n_1488), .Y (n_1470));
NAND2X1 g39814(.A (u8_mem_b2_b_50 ), .B (n_2366), .Y (n_2244));
AOI22X1 g37645(.A0 (n_6933), .A1 (n_1835), .B0 (n_6915), .B1(n_1760), .Y (n_1718));
NAND2X1 g39815(.A (n_2344), .B (in_slt_421), .Y (n_1901));
NAND2X1 g39816(.A (n_3259), .B (u5_mem_b0_b_103 ), .Y (n_12855));
INVX1 g41232(.A (n_2463), .Y (n_1404));
NAND2X1 g39817(.A (u7_mem_b1_b_64 ), .B (n_3522), .Y (n_2943));
INVX8 g41231(.A (n_1052), .Y (n_2463));
NOR2X1 g35353(.A (i3_status), .B (i3_status_1022), .Y (n_7032));
NOR2X1 g41230(.A (u11_rp_b0_b ), .B (u11_wp_b1_b ), .Y (n_916));
NOR2X1 g41237(.A (n_63), .B (n_600), .Y (n_839));
OAI21X1 g33000(.A0 (n_7269), .A1 (n_6998), .B0 (n_12609), .Y(n_9815));
NAND2X1 g39673(.A (n_996), .B (wb_addr_i_b4_b), .Y (n_1216));
INVX2 g41235(.A (n_839), .Y (n_1052));
AOI22X1 g37926(.A0 (u9_din_tmp_51), .A1 (n_2368), .B0 (in_slt_408),.B1 (n_4624), .Y (n_2633));
NAND2X1 g39674(.A (u7_mem_b2_b_57 ), .B (n_12650), .Y (n_4148));
NAND2X1 g39675(.A (u4_mem_b1_b_78 ), .B (n_12259), .Y (n_4147));
AOI21X1 g38563(.A0 (u8_mem_b1_b_67 ), .A1 (n_4502), .B0 (n_2068), .Y(n_4274));
NOR2X1 g35355(.A (i6_status), .B (i6_status_1042), .Y (n_7157));
AOI21X1 g38562(.A0 (u8_mem_b1_b_68 ), .A1 (n_4387), .B0 (n_2069), .Y(n_4275));
NOR2X1 g39677(.A (u11_mem_b2_b ), .B (n_1214), .Y (n_1215));
AOI21X1 g38561(.A0 (u3_mem_b1_b_73 ), .A1 (n_5157), .B0 (n_2757), .Y(n_4867));
AOI21X1 g38560(.A0 (u5_mem_b2_b_47 ), .A1 (n_4378), .B0 (n_1932), .Y(n_4276));
NAND2X1 g39601(.A (u5_mem_b1_b_82 ), .B (n_3239), .Y (n_3069));
AOI21X1 g38567(.A0 (u3_mem_b1_b_78 ), .A1 (n_5148), .B0 (n_2819), .Y(n_4864));
AOI21X1 g38566(.A0 (u3_mem_b1_b_76 ), .A1 (n_5148), .B0 (n_2813), .Y(n_4865));
INVX2 g35046(.A (n_7414), .Y (n_8333));
AOI21X1 g38565(.A0 (u8_mem_b2_b_38 ), .A1 (n_4491), .B0 (n_1979), .Y(n_4273));
INVX2 g35040(.A (n_7414), .Y (n_9349));
AOI21X1 g38564(.A0 (u3_mem_b1_b_75 ), .A1 (n_5157), .B0 (n_2839), .Y(n_4866));
NAND2X1 g39600(.A (n_12204), .B (u6_mem_b0_b_117 ), .Y (n_3070));
INVX1 g42027(.A (u11_mem_b2_b_117 ), .Y (n_190));
INVX1 g42025(.A (u10_mem_b1_b_140 ), .Y (n_87));
INVX1 g42024(.A (n_4708), .Y (n_872));
INVX1 g42022(.A (ic0_cfg_1029), .Y (n_410));
INVX1 g42021(.A (n_410), .Y (n_4699));
INVX1 g42020(.A (u9_mem_b3_b_76 ), .Y (n_5294));
INVX1 g42029(.A (u10_mem_b0_b_157 ), .Y (n_5945));
INVX8 g35223(.A (n_7976), .Y (n_7490));
AOI21X1 g35954(.A0 (n_6972), .A1 (n_862), .B0 (n_5791), .Y (n_6974));
AOI21X1 g35957(.A0 (n_6972), .A1 (oc1_cfg_980), .B0 (n_5763), .Y(n_6969));
AOI21X1 g35956(.A0 (n_6972), .A1 (n_8565), .B0 (n_5765), .Y (n_6971));
OAI21X1 g35951(.A0 (n_5567), .A1 (n_7063), .B0 (n_5899), .Y (n_6975));
OAI21X1 g35953(.A0 (n_6082), .A1 (n_11934), .B0 (n_6791), .Y(n_7175));
OAI21X1 g35952(.A0 (n_5572), .A1 (n_7063), .B0 (n_6261), .Y (n_7052));
NAND2X1 g39216(.A (n_12840), .B (u4_mem_b0_b_111 ), .Y (n_3362));
NAND2X1 g39217(.A (u8_mem_b1_b_73 ), .B (n_12295), .Y (n_11458));
INVX1 g39214(.A (n_4764), .Y (n_3363));
NAND2X1 g39215(.A (in_slt_414), .B (n_2368), .Y (n_4764));
AOI21X1 g35959(.A0 (n_6972), .A1 (oc0_cfg_966), .B0 (n_5785), .Y(n_6967));
AOI21X1 g35958(.A0 (n_6972), .A1 (oc0_cfg_965), .B0 (n_5787), .Y(n_6968));
NOR2X1 g39210(.A (n_3089), .B (n_2712), .Y (n_3370));
NAND2X1 g39211(.A (u4_mem_b2_b_48 ), .B (n_12087), .Y (n_3367));
NAND2X1 g36914(.A (n_1672), .B (n_1671), .Y (n_4032));
INVX4 g45968_dup(.A (n_12735), .Y (n_12826));
OAI21X1 g33408(.A0 (n_3867), .A1 (n_8894), .B0 (n_8154), .Y (n_8468));
NAND2X1 g34794(.A (u7_mem_b3_b_142 ), .B (n_7651), .Y (n_7639));
NAND2X1 g34795(.A (u7_mem_b3_b_143 ), .B (n_7651), .Y (n_7638));
NAND2X1 g34796(.A (u7_mem_b3_b_144 ), .B (n_7651), .Y (n_7637));
NAND2X1 g34790(.A (u7_mem_b3_b_139 ), .B (n_7651), .Y (n_7643));
NAND2X1 g34791(.A (u7_mem_b3_b_140 ), .B (n_7651), .Y (n_7642));
NAND2X1 g34792(.A (u7_mem_b3_b_122 ), .B (n_7651), .Y (n_7641));
NAND2X1 g34793(.A (u7_mem_b3_b_141 ), .B (n_7651), .Y (n_7640));
NAND2X1 g38826(.A (u8_mem_b3_b_124 ), .B (n_2468), .Y (n_2453));
NAND2X1 g34798(.A (u7_mem_b3_b_146 ), .B (n_7651), .Y (n_7635));
NAND2X1 g34799(.A (u7_mem_b3_b_147 ), .B (n_7651), .Y (n_7634));
NAND2X1 g39581(.A (n_12204), .B (u6_mem_b0_b_102 ), .Y (n_11697));
NAND2X1 g38827(.A (u6_mem_b3_b_133 ), .B (n_12622), .Y (n_2452));
NOR2X1 g34887(.A (o3_status), .B (o3_status_962), .Y (n_7166));
NAND2X1 g34570(.A (u5_mem_b3_b_144 ), .B (n_7870), .Y (n_7856));
NAND2X1 g34571(.A (u5_mem_b3_b_145 ), .B (n_7870), .Y (n_7855));
NAND2X1 g34572(.A (u5_mem_b3_b_146 ), .B (n_7870), .Y (n_7854));
NAND2X1 g34573(.A (u5_mem_b3_b_147 ), .B (n_7870), .Y (n_7853));
NAND2X1 g34574(.A (u5_mem_b3_b_148 ), .B (n_7870), .Y (n_7852));
NAND2X1 g34575(.A (u5_mem_b3_b_149 ), .B (n_7870), .Y (n_7851));
NAND2X1 g34576(.A (u5_mem_b3_b_150 ), .B (n_7870), .Y (n_7850));
NAND2X1 g34577(.A (u5_mem_b3_b_123 ), .B (n_7870), .Y (n_7849));
NAND2X1 g34578(.A (u5_mem_b3_b_151 ), .B (n_7870), .Y (n_7848));
NAND2X1 g34579(.A (u5_mem_b3_b_152 ), .B (n_7870), .Y (n_7847));
INVX1 g41824(.A (u10_mem_b1_b_144 ), .Y (n_1676));
INVX4 g41822(.A (n_2567), .Y (n_6152));
INVX4 g41823(.A (n_610), .Y (n_2567));
NAND2X1 g38948(.A (u6_mem_b3_b_126 ), .B (n_12622), .Y (n_2398));
INVX1 g43088(.A (u10_mem_b3_b_81 ), .Y (n_5512));
INVX1 g43089(.A (u10_mem_b0_b_177 ), .Y (n_1238));
INVX1 g43086(.A (wb_ack_o), .Y (n_303));
NAND2X1 g41022(.A (n_808), .B (n_4711), .Y (n_7080));
INVX1 g43084(.A (u11_mem_b2_b_90 ), .Y (n_6445));
INVX1 g43083(.A (u9_mem_b2_b_91 ), .Y (n_6931));
INVX1 g43081(.A (u9_mem_b1_b_146 ), .Y (n_1723));
AND2X1 g34881(.A (u15_valid_r), .B (n_11827), .Y (n_9710));
CLKBUFX1 g45613(.A (n_12281), .Y (n_12280));
AOI21X1 g38146(.A0 (u4_mem_b2_b_41 ), .A1 (n_4439), .B0 (n_2170), .Y(n_4438));
NAND2X1 g39763(.A (n_4560), .B (in_slt_456), .Y (n_5304));
AOI22X1 g37635(.A0 (n_340), .A1 (n_1859), .B0 (n_5372), .B1 (n_1760),.Y (n_1735));
NAND2X1 g39766(.A (n_3252), .B (u7_mem_b0_b_121 ), .Y (n_2970));
INVX1 g42840(.A (n_626), .Y (n_6838));
INVX1 g42845(.A (u10_mem_b1_b_128 ), .Y (n_6476));
INVX1 g42847(.A (u11_mem_b2_b_96 ), .Y (n_5969));
INVX1 g42846(.A (u9_mem_b1_b_131 ), .Y (n_6534));
NAND2X1 g37171(.A (n_2516), .B (n_2197), .Y (n_5987));
NAND2X1 g37170(.A (n_2519), .B (n_2261), .Y (n_6011));
AOI21X1 g38301(.A0 (u5_mem_b1_b_68 ), .A1 (n_5048), .B0 (n_2731), .Y(n_5010));
NAND2X1 g37172(.A (n_3898), .B (n_2326), .Y (n_6453));
NAND2X1 g37175(.A (n_3896), .B (n_2472), .Y (n_6497));
NAND2X1 g37174(.A (n_3899), .B (n_2270), .Y (n_6589));
AOI21X1 g38304(.A0 (u7_mem_b1_b_90 ), .A1 (n_5118), .B0 (n_2837), .Y(n_5009));
NAND2X1 g37179(.A (n_4566), .B (n_2296), .Y (n_6544));
NAND2X1 g37178(.A (n_4567), .B (n_2251), .Y (n_6442));
AOI21X1 g38309(.A0 (u5_mem_b2_b_42 ), .A1 (n_4378), .B0 (n_1933), .Y(n_4374));
AOI21X1 g38308(.A0 (u6_mem_b1_b_84 ), .A1 (n_5019), .B0 (n_2820), .Y(n_5008));
NAND2X1 g36559(.A (n_5818), .B (n_6773), .Y (n_5819));
NAND2X1 g36554(.A (n_6202), .B (n_6201), .Y (n_6203));
NAND2X1 g36556(.A (n_6228), .B (n_6201), .Y (n_6200));
NAND2X1 g36557(.A (n_12514), .B (n_6201), .Y (n_6199));
NAND2X1 g36552(.A (n_6204), .B (n_6773), .Y (n_6205));
INVX1 g42908(.A (oc3_cfg_995), .Y (n_319));
INVX1 g42909(.A (u10_mem_b0_b_172 ), .Y (n_1242));
INVX1 g42904(.A (oc3_cfg_997), .Y (n_571));
INVX4 g45625(.A (n_12304), .Y (n_12303));
INVX1 g42906(.A (u9_mem_b1_b_123 ), .Y (n_6945));
INVX1 g42907(.A (u10_mem_b0_b_152 ), .Y (n_6339));
INVX1 g42900(.A (u10_mem_b1_b_149 ), .Y (n_162));
INVX1 g42902(.A (u10_mem_b0_b_171 ), .Y (n_2557));
INVX4 g45623(.A (n_12303), .Y (n_12295));
NAND2X1 g39764(.A (n_2325), .B (in_slt_445), .Y (n_2296));
INVX1 g35133(.A (n_7408), .Y (n_9264));
NAND2X1 g38918(.A (u7_mem_b3_b_142 ), .B (n_1546), .Y (n_1347));
NAND2X1 g40995(.A (n_8526), .B (n_924), .Y (n_9591));
AOI22X1 g37795(.A0 (n_2558), .A1 (n_6335), .B0 (n_6623), .B1(n_2544), .Y (n_1646));
NAND2X1 g37794(.A (n_4134), .B (n_3422), .Y (n_5213));
NAND2X1 g37797(.A (n_2429), .B (n_2908), .Y (n_12055));
AOI22X1 g37791(.A0 (n_2558), .A1 (n_6337), .B0 (n_6572), .B1(n_1316), .Y (n_1236));
AOI22X1 g37790(.A0 (n_5978), .A1 (n_1575), .B0 (n_6026), .B1(n_1831), .Y (n_1652));
AOI22X1 g37793(.A0 (n_129), .A1 (n_1575), .B0 (n_5580), .B1 (n_1831),.Y (n_1648));
AOI22X1 g37792(.A0 (n_1756), .A1 (n_334), .B0 (n_1650), .B1 (n_1643),.Y (n_1651));
AOI22X1 g37799(.A0 (n_6411), .A1 (n_1839), .B0 (n_6569), .B1(n_1316), .Y (n_1640));
AOI22X1 g37798(.A0 (n_288), .A1 (n_1575), .B0 (n_5582), .B1 (n_1831),.Y (n_1642));
OAI21X1 g33085(.A0 (n_7172), .A1 (n_6975), .B0 (n_10483), .Y(n_11631));
OAI21X1 g33084(.A0 (n_7276), .A1 (n_6976), .B0 (n_10483), .Y(n_11639));
OAI21X1 g33087(.A0 (n_7275), .A1 (n_7177), .B0 (n_9885), .Y(n_11984));
OAI21X1 g33086(.A0 (n_7114), .A1 (n_7052), .B0 (n_10483), .Y(n_11641));
OAI21X1 g33081(.A0 (n_7207), .A1 (n_7054), .B0 (n_10483), .Y(n_11635));
OAI21X1 g33080(.A0 (n_7208), .A1 (n_7055), .B0 (n_10481), .Y(n_12016));
OAI21X1 g33083(.A0 (n_7204), .A1 (n_6977), .B0 (n_10483), .Y(n_11637));
OAI21X1 g33082(.A0 (n_7205), .A1 (n_7053), .B0 (n_10483), .Y(n_11992));
MX2X1 g33089(.A (n_392), .B (wb_din), .S0 (n_8643), .Y (n_8655));
OAI21X1 g33088(.A0 (n_9711), .A1 (u15_rdd2), .B0 (n_716), .Y(n_9796));
NOR2X1 g41209(.A (n_8565), .B (n_942), .Y (n_9768));
OAI21X1 g31029(.A0 (n_5281), .A1 (n_10820), .B0 (n_10382), .Y(n_10888));
OAI21X1 g31028(.A0 (n_5327), .A1 (n_10880), .B0 (n_10383), .Y(n_10890));
AOI21X1 g31799(.A0 (n_10983), .A1 (n_10617), .B0 (n_10614), .Y(n_10984));
AOI21X1 g31798(.A0 (n_4068), .A1 (n_9481), .B0 (n_9495), .Y (n_9482));
OAI21X1 g31025(.A0 (n_5323), .A1 (n_10820), .B0 (n_10387), .Y(n_10894));
AOI21X1 g31796(.A0 (n_1411), .A1 (n_1845), .B0 (n_11892), .Y(n_9963));
OAI21X1 g31027(.A0 (n_5329), .A1 (n_10880), .B0 (n_10384), .Y(n_10892));
OAI21X1 g31026(.A0 (n_5332), .A1 (n_10820), .B0 (n_10386), .Y(n_10893));
OAI21X1 g31021(.A0 (n_5415), .A1 (n_10450), .B0 (n_9992), .Y(n_10677));
OAI21X1 g31020(.A0 (n_5416), .A1 (n_10880), .B0 (n_10392), .Y(n_10898));
AOI21X1 g31791(.A0 (n_10988), .A1 (n_9876), .B0 (n_10633), .Y(n_10989));
OAI21X1 g31022(.A0 (n_5414), .A1 (n_10880), .B0 (n_10390), .Y(n_10897));
INVX1 g42447(.A (u11_mem_b3_b_59 ), .Y (n_6417));
INVX1 g40873(.A (n_1430), .Y (n_2713));
NAND2X1 g41018(.A (n_8197), .B (n_804), .Y (n_9585));
NAND3X1 g33337(.A (n_1873), .B (n_7048), .C (n_7758), .Y (n_8177));
NAND4X1 g33336(.A (n_5618), .B (n_1806), .C (n_7505), .D (n_1256), .Y(n_9450));
NOR2X1 g33335(.A (n_11529), .B (n_8665), .Y (n_9569));
INVX1 g33334(.A (n_9569), .Y (n_9668));
INVX1 g33333(.A (n_9668), .Y (n_9705));
INVX4 g33332(.A (n_9705), .Y (n_9876));
INVX4 g41011(.A (n_1221), .Y (n_1835));
NAND2X1 g41010(.A (n_590), .B (oc5_cfg_1016), .Y (n_928));
AOI22X1 g37934(.A0 (n_2502), .A1 (n_2507), .B0 (n_2506), .B1(n_1859), .Y (n_2508));
BUFX3 g40870(.A (n_1226), .Y (n_5118));
AOI22X1 g37937(.A0 (n_236), .A1 (n_1575), .B0 (n_5502), .B1 (n_1831),.Y (n_1855));
MX2X1 g31249(.A (n_6403), .B (n_6402), .S0 (n_10308), .Y (n_10173));
MX2X1 g31241(.A (n_5967), .B (n_5966), .S0 (n_10315), .Y (n_10179));
MX2X1 g31240(.A (n_6443), .B (n_6441), .S0 (n_10513), .Y (n_10452));
MX2X1 g31243(.A (n_6659), .B (n_6658), .S0 (n_9818), .Y (n_10828));
MX2X1 g31242(.A (n_6557), .B (n_6556), .S0 (n_10839), .Y (n_10829));
MX2X1 g31245(.A (n_6626), .B (n_6625), .S0 (n_9818), .Y (n_10827));
MX2X1 g31244(.A (n_6038), .B (n_6037), .S0 (n_10315), .Y (n_10178));
MX2X1 g31247(.A (n_6869), .B (n_6868), .S0 (n_10308), .Y (n_10176));
XOR2X1 g31246(.A (n_610), .B (n_9908), .Y (n_10825));
NAND2X1 g39681(.A (u6_mem_b2_b_43 ), .B (n_2285), .Y (n_2264));
NAND2X1 g39683(.A (n_2302), .B (in_slt_423), .Y (n_2261));
NOR2X1 g39685(.A (n_3486), .B (n_2712), .Y (n_2810));
OAI21X1 g33563(.A0 (n_4416), .A1 (n_9326), .B0 (n_7994), .Y (n_8273));
NOR2X1 g39686(.A (n_3332), .B (n_2748), .Y (n_3022));
NAND2X1 g39689(.A (n_2513), .B (in_slt_445), .Y (n_2197));
NAND2X1 g39688(.A (u11_din_tmp_50), .B (n_4560), .Y (n_3020));
NAND2X1 g38796(.A (u4_mem_b3_b_135 ), .B (n_12744), .Y (n_11651));
NAND2X1 g38797(.A (u3_mem_b3_b_145 ), .B (n_2463), .Y (n_2459));
NOR2X1 g38798(.A (n_421), .B (wb_addr_i_b30_b), .Y (n_1262));
NAND2X1 g38799(.A (n_605), .B (n_1142), .Y (n_3942));
NOR2X1 g41145(.A (n_4703), .B (n_872), .Y (n_8847));
CLKBUFX3 g40699(.A (n_1178), .Y (n_2362));
NOR2X1 g41412(.A (u13_ints_r_b18_b ), .B (n_611), .Y (n_612));
NAND2X1 g37562(.A (n_5645), .B (n_4178), .Y (n_5235));
INVX2 g40690(.A (n_933), .Y (n_1180));
INVX1 g40691(.A (n_1180), .Y (n_2045));
NAND2X2 g40696(.A (u8_wp_b0_b ), .B (n_178), .Y (n_933));
OR2X1 g41411(.A (n_454), .B (n_418), .Y (n_847));
INVX2 g41141(.A (n_1149), .Y (n_1411));
CLKBUFX1 g45822(.A (n_12534), .Y (n_12535));
AND2X1 g45823(.A (n_257), .B (n_925), .Y (n_12534));
OAI21X1 g45820(.A0 (n_4601), .A1 (n_4600), .B0 (n_12536), .Y(n_12537));
AND2X1 g45821(.A (n_634), .B (n_12535), .Y (n_12536));
NAND2X1 g41143(.A (u6_rp_b2_b ), .B (n_11579), .Y (n_781));
NAND3X1 g45824(.A (n_6316), .B (n_12535), .C (n_6163), .Y (n_12538));
INVX2 g41414(.A (n_736), .Y (n_1831));
AOI21X1 g35564(.A0 (n_6312), .A1 (n_6137), .B0 (n_7324), .Y (n_7279));
NOR2X1 g30045(.A (n_12585), .B (n_11526), .Y (n_11181));
NOR2X1 g30046(.A (n_11142), .B (n_5839), .Y (n_11180));
NOR2X1 g30047(.A (n_1870), .B (n_11520), .Y (n_11179));
NAND2X1 g35560(.A (n_6045), .B (n_5225), .Y (n_7025));
NAND2X1 g35561(.A (n_6045), .B (n_6044), .Y (n_7022));
NAND2X1 g35562(.A (n_6045), .B (n_6042), .Y (n_6043));
AND2X1 g35563(.A (n_5226), .B (n_2608), .Y (n_6041));
NOR2X1 g30048(.A (n_5825), .B (n_11522), .Y (n_11178));
NAND3X1 g30049(.A (n_9702), .B (n_9525), .C (n_9616), .Y (n_9850));
INVX1 g40875(.A (n_1430), .Y (n_2836));
NAND2X1 g37543(.A (n_553), .B (in_slt_742), .Y (n_1023));
BUFX3 g40832(.A (n_867), .Y (n_4378));
INVX1 g34962(.A (n_7428), .Y (n_9165));
INVX4 g39105(.A (n_1185), .Y (n_5272));
INVX1 g34966(.A (n_7428), .Y (n_9139));
NOR2X1 g39022(.A (n_3332), .B (n_2804), .Y (n_3507));
BUFX3 g34969(.A (o7_we), .Y (n_7428));
NAND2X1 g31718(.A (n_5526), .B (n_10385), .Y (n_10355));
OAI21X1 g35876(.A0 (n_5714), .A1 (n_6995), .B0 (n_5878), .Y (n_7162));
OAI21X1 g35877(.A0 (n_5562), .A1 (n_6995), .B0 (n_5877), .Y (n_6996));
OAI21X1 g35874(.A0 (n_5564), .A1 (n_7115), .B0 (n_5883), .Y (n_6993));
OAI21X1 g35873(.A0 (n_5716), .A1 (n_7115), .B0 (n_5885), .Y (n_7102));
NAND2X1 g37162(.A (n_4584), .B (n_2940), .Y (n_6913));
AOI21X1 g35654(.A0 (n_5909), .A1 (n_5790), .B0 (n_7120), .Y (n_7119));
AOI21X1 g38315(.A0 (u5_mem_b2_b_48 ), .A1 (n_4370), .B0 (n_2055), .Y(n_4367));
AOI21X1 g38316(.A0 (u7_mem_b2_b_33 ), .A1 (n_4509), .B0 (n_2035), .Y(n_4366));
NAND2X1 g34703(.A (u3_mem_b1_b_74 ), .B (n_8101), .Y (n_7725));
AOI21X1 g38317(.A0 (u5_mem_b2_b_49 ), .A1 (n_4370), .B0 (n_1954), .Y(n_4365));
AOI21X1 g38310(.A0 (u5_mem_b2_b_43 ), .A1 (n_4370), .B0 (n_2198), .Y(n_4373));
NAND2X1 g34701(.A (u8_mem_b1_b_66 ), .B (n_7976), .Y (n_7726));
AOI21X1 g38311(.A0 (u5_mem_b2_b_44 ), .A1 (n_4378), .B0 (n_2167), .Y(n_4372));
NOR2X1 g34700(.A (o8_status_1002), .B (n_5825), .Y (n_9483));
AND2X1 g40937(.A (n_708), .B (u10_wp_b2_b ), .Y (n_931));
AOI21X1 g38312(.A0 (u5_mem_b2_b_45 ), .A1 (n_4370), .B0 (n_2042), .Y(n_4371));
NAND2X1 g34871(.A (u8_mem_b2_b_57 ), .B (n_7976), .Y (n_7563));
AOI21X1 g38313(.A0 (u5_mem_b2_b_46 ), .A1 (n_4370), .B0 (n_2226), .Y(n_4369));
NAND3X1 g34706(.A (n_4703), .B (n_4708), .C (n_865), .Y (n_1887));
OR2X1 g34705(.A (i3_status), .B (n_7383), .Y (n_7384));
AOI21X1 g35677(.A0 (n_1000), .A1 (n_1214), .B0 (i6_re), .Y (n_6750));
NAND2X1 g34704(.A (n_7385), .B (n_7383), .Y (n_7532));
MX2X1 g38648(.A (u5_mem_b0_b_102 ), .B (wb_din_672), .S0 (n_3720), .Y(n_3735));
OAI21X1 g33535(.A0 (n_4297), .A1 (n_8333), .B0 (n_8022), .Y (n_8306));
OAI21X1 g33534(.A0 (n_4446), .A1 (n_9336), .B0 (n_8023), .Y (n_8308));
OAI21X1 g33537(.A0 (n_4444), .A1 (n_8333), .B0 (n_8020), .Y (n_8304));
OAI21X1 g33536(.A0 (n_4445), .A1 (n_8318), .B0 (n_8021), .Y (n_8305));
OAI21X1 g33531(.A0 (n_4449), .A1 (n_8333), .B0 (n_8026), .Y (n_8311));
OAI21X1 g33530(.A0 (n_4450), .A1 (n_9326), .B0 (n_8027), .Y (n_8313));
OAI21X1 g33533(.A0 (n_4447), .A1 (n_9336), .B0 (n_8024), .Y (n_8309));
OAI21X1 g33532(.A0 (n_4448), .A1 (n_8333), .B0 (n_8025), .Y (n_8310));
OAI21X1 g33539(.A0 (n_4442), .A1 (n_8333), .B0 (n_8018), .Y (n_8302));
OAI21X1 g33538(.A0 (n_4295), .A1 (n_9349), .B0 (n_8019), .Y (n_8303));
NAND2X1 g34466(.A (u4_mem_b3_b_125 ), .B (n_7984), .Y (n_7955));
OR2X1 g46001(.A (n_485), .B (n_422), .Y (n_12801));
INVX8 g46003(.A (n_12401), .Y (n_12823));
NAND2X1 g37548(.A (n_974), .B (in_slt_742), .Y (n_1259));
NAND2X1 g37549(.A (n_811), .B (in_slt_742), .Y (n_1289));
OR2X1 g46002(.A (n_524), .B (n_447), .Y (n_12803));
INVX1 g37092(.A (n_6176), .Y (n_5676));
NAND4X1 g37093(.A (n_3183), .B (n_1487), .C (n_3126), .D (n_1512), .Y(n_6176));
NAND4X1 g37090(.A (n_11451), .B (n_11452), .C (n_2353), .D (n_2457),.Y (n_5813));
NAND4X1 g37091(.A (n_3469), .B (n_2894), .C (n_3227), .D (n_2392), .Y(n_6165));
INVX1 g37096(.A (n_6182), .Y (n_5675));
INVX1 g37094(.A (n_5811), .Y (n_5532));
NAND4X1 g37095(.A (n_11459), .B (n_11460), .C (n_2299), .D (n_2373),.Y (n_5811));
OAI21X1 g33658(.A0 (n_4300), .A1 (n_9286), .B0 (n_7882), .Y (n_9247));
OAI21X1 g33659(.A0 (n_4301), .A1 (n_9286), .B0 (n_7881), .Y (n_9246));
CLKBUFX1 g46007(.A (n_12848), .Y (n_12847));
OAI21X1 g33650(.A0 (n_4364), .A1 (n_9307), .B0 (n_7890), .Y (n_9257));
OAI21X1 g33651(.A0 (n_4289), .A1 (n_9286), .B0 (n_7889), .Y (n_9256));
OAI21X1 g33652(.A0 (n_4363), .A1 (n_9264), .B0 (n_7888), .Y (n_9255));
OAI21X1 g33653(.A0 (n_4362), .A1 (n_9264), .B0 (n_7887), .Y (n_9254));
OAI21X1 g33654(.A0 (n_4361), .A1 (n_9235), .B0 (n_7886), .Y (n_9253));
OAI21X1 g33655(.A0 (n_4360), .A1 (n_9202), .B0 (n_7885), .Y (n_9252));
OAI21X1 g33657(.A0 (n_4357), .A1 (n_9264), .B0 (n_7883), .Y (n_9249));
AOI21X1 g38516(.A0 (u7_mem_b3_b_142 ), .A1 (n_4961), .B0 (n_3076), .Y(n_4883));
INVX1 g37325(.A (n_4728), .Y (n_5275));
AOI21X1 g38514(.A0 (u7_mem_b3_b_127 ), .A1 (n_4961), .B0 (n_3381), .Y(n_4885));
AOI21X1 g38515(.A0 (u7_mem_b3_b_122 ), .A1 (n_4961), .B0 (n_3409), .Y(n_4884));
AOI22X1 g37320(.A0 (n_5272), .A1 (u13_intm_r_b0_b ), .B0 (n_5277), .B1(crac_din), .Y (n_5278));
AOI22X1 g37321(.A0 (n_5591), .A1 (n_11772), .B0 (n_6972), .B1(n_997), .Y (n_4733));
AOI21X1 g38510(.A0 (u7_mem_b3_b_133 ), .A1 (n_5145), .B0 (n_3520), .Y(n_4887));
AOI22X1 g37323(.A0 (n_5272), .A1 (u13_intm_r_b1_b ), .B0 (n_5277), .B1(crac_din_692), .Y (n_5276));
AOI22X1 g37898(.A0 (n_2325), .A1 (in_slt_458), .B0 (n_2513), .B1(in_slt_446), .Y (n_5413));
AOI22X1 g37899(.A0 (n_2325), .A1 (in_slt_459), .B0 (n_2513), .B1(in_slt_447), .Y (n_5410));
INVX1 g37328(.A (n_3991), .Y (n_4725));
AOI22X1 g37329(.A0 (n_5277), .A1 (crac_out_866), .B0 (n_6972), .B1(n_8550), .Y (n_3991));
AOI21X1 g38518(.A0 (u7_mem_b3_b_146 ), .A1 (n_5145), .B0 (n_2976), .Y(n_4881));
AOI21X1 g38519(.A0 (u5_mem_b2_b_58 ), .A1 (n_4370), .B0 (n_2172), .Y(n_4301));
MX2X1 g36089(.A (n_6492), .B (n_6444), .S0 (n_995), .Y (n_6493));
INVX1 g45611(.A (n_12280), .Y (n_12278));
NAND2X1 g38868(.A (u4_mem_b3_b_148 ), .B (n_3556), .Y (n_3538));
NAND2X1 g34639(.A (u6_mem_b2_b_43 ), .B (n_7758), .Y (n_7786));
NAND2X1 g38862(.A (u5_mem_b3_b_124 ), .B (n_3543), .Y (n_2438));
INVX4 g40930(.A (n_931), .Y (n_1162));
NAND2X1 g38863(.A (u5_mem_b3_b_125 ), .B (n_1543), .Y (n_1338));
OAI21X1 g33486(.A0 (n_5129), .A1 (n_8372), .B0 (n_8085), .Y (n_8367));
NAND2X1 g38860(.A (u5_mem_b3_b_123 ), .B (n_1543), .Y (n_1335));
AOI21X1 g37301(.A0 (n_5302), .A1 (n_5371), .B0 (n_3947), .Y (n_5303));
NAND2X1 g32703(.A (n_79), .B (n_10617), .Y (n_10619));
NAND2X1 g38867(.A (u4_mem_b3_b_137 ), .B (n_3546), .Y (n_3539));
NAND2X1 g38864(.A (u3_mem_b3_b_148 ), .B (n_2463), .Y (n_2437));
NAND2X1 g38865(.A (u5_mem_b3_b_126 ), .B (n_1543), .Y (n_1337));
BUFX3 g41466(.A (n_4996), .Y (n_5000));
NOR2X1 g41464(.A (u13_ints_r_b22_b ), .B (n_739), .Y (n_740));
AOI21X1 g38184(.A0 (u7_mem_b2_b_38 ), .A1 (n_4540), .B0 (n_2087), .Y(n_4406));
MX2X1 g36055(.A (n_6551), .B (n_6618), .S0 (n_4783), .Y (n_6552));
MX2X1 g36054(.A (n_6521), .B (n_6554), .S0 (n_6649), .Y (n_6555));
MX2X1 g36057(.A (n_6548), .B (n_6547), .S0 (n_995), .Y (n_6549));
MX2X1 g36056(.A (n_6899), .B (n_6886), .S0 (n_6908), .Y (n_6887));
MX2X1 g36051(.A (n_6891), .B (n_6890), .S0 (n_6908), .Y (n_6892));
MX2X1 g36050(.A (n_5998), .B (n_5997), .S0 (n_5341), .Y (n_5999));
MX2X1 g36053(.A (n_6544), .B (n_6556), .S0 (n_6649), .Y (n_6557));
MX2X1 g36052(.A (n_6888), .B (n_6891), .S0 (n_930), .Y (n_6889));
MX2X1 g36059(.A (n_6884), .B (n_6883), .S0 (n_4783), .Y (n_6885));
MX2X1 g36058(.A (n_6545), .B (n_6544), .S0 (n_6502), .Y (n_6546));
INVX4 g42042(.A (n_3559), .Y (n_5772));
INVX4 g42045(.A (n_6091), .Y (n_3559));
INVX1 g42047(.A (u10_mem_b2_b_96 ), .Y (n_6018));
INVX1 g42046(.A (u9_mem_b3_b_78 ), .Y (n_5343));
NOR2X1 g40308(.A (n_945), .B (n_2702), .Y (n_1971));
NAND2X1 g39238(.A (u6_mem_b1_b_72 ), .B (n_4253), .Y (n_11700));
NOR2X1 g39239(.A (n_4961), .B (n_2792), .Y (n_3535));
INVX1 g40759(.A (n_1174), .Y (n_2216));
BUFX3 g40758(.A (n_938), .Y (n_4509));
MX2X1 g35979(.A (n_6028), .B (n_6008), .S0 (n_931), .Y (n_6029));
MX2X1 g35978(.A (n_6030), .B (n_6011), .S0 (n_931), .Y (n_6031));
MX2X1 g35977(.A (n_6033), .B (n_6014), .S0 (n_5341), .Y (n_6034));
MX2X1 g35976(.A (n_6660), .B (n_6586), .S0 (n_5341), .Y (n_6661));
MX2X1 g35975(.A (n_6662), .B (n_6589), .S0 (n_5341), .Y (n_6663));
MX2X1 g35974(.A (n_6664), .B (n_6592), .S0 (n_5341), .Y (n_6665));
MX2X1 g35973(.A (n_6666), .B (n_6596), .S0 (n_5341), .Y (n_6667));
MX2X1 g35972(.A (n_6668), .B (n_6599), .S0 (n_931), .Y (n_6669));
MX2X1 g35970(.A (n_5983), .B (n_6035), .S0 (n_6649), .Y (n_6036));
CLKBUFX1 g42372(.A (u10_wp_b1_b ), .Y (n_5420));
NOR2X1 g40306(.A (n_2477), .B (n_2772), .Y (n_1973));
NAND2X1 g34633(.A (u6_mem_b2_b_38 ), .B (n_7758), .Y (n_7792));
NOR2X1 g40266(.A (n_2020), .B (n_2720), .Y (n_2000));
NOR2X1 g40301(.A (n_2099), .B (n_2735), .Y (n_1976));
NOR2X1 g40265(.A (n_2763), .B (n_1985), .Y (n_1871));
INVX1 g42639(.A (oc4_int_set_716), .Y (n_463));
INVX1 g41805(.A (u4_wp_b2_b ), .Y (n_95));
NAND2X1 g34778(.A (u7_mem_b2_b_35 ), .B (n_7651), .Y (n_7656));
NAND2X1 g34779(.A (u7_mem_b2_b_36 ), .B (n_7651), .Y (n_7655));
NAND2X1 g34776(.A (u7_mem_b2_b_33 ), .B (n_7651), .Y (n_7658));
NAND2X1 g34774(.A (u7_mem_b2_b_31 ), .B (n_7651), .Y (n_7660));
NAND2X1 g34775(.A (u7_mem_b2_b_32 ), .B (n_7651), .Y (n_7659));
NAND2X1 g34772(.A (u8_mem_b2_b_52 ), .B (n_7976), .Y (n_7662));
NAND2X1 g34773(.A (u7_mem_b2_b_59 ), .B (n_7651), .Y (n_7661));
NAND2X1 g34770(.A (u7_mem_b2_b_30 ), .B (n_7651), .Y (n_7664));
NAND2X1 g34771(.A (u7_mem_b2_b_58 ), .B (n_7651), .Y (n_7663));
NOR2X1 g39010(.A (n_2801), .B (n_1488), .Y (n_1503));
INVX2 g40645(.A (wb_din_688), .Y (n_2767));
NOR2X1 g39991(.A (n_2763), .B (n_2067), .Y (n_2214));
BUFX3 g41696(.A (n_4961), .Y (n_5145));
INVX1 g41808(.A (u11_mem_b1_b_122 ), .Y (n_6490));
INVX1 g41809(.A (u11_mem_b2_b_97 ), .Y (n_6479));
NAND2X1 g34518(.A (u5_mem_b1_b_65 ), .B (n_7870), .Y (n_7910));
NAND2X1 g34519(.A (u5_mem_b1_b_66 ), .B (n_7870), .Y (n_7909));
NAND2X1 g34512(.A (u5_mem_b1_b_61 ), .B (n_7870), .Y (n_7916));
NAND2X1 g34513(.A (u5_mem_b1_b_89 ), .B (n_7870), .Y (n_7915));
NAND2X1 g34510(.A (u5_mem_b1_b_87 ), .B (n_7870), .Y (n_7918));
NAND2X1 g34511(.A (u5_mem_b1_b_88 ), .B (n_7870), .Y (n_7917));
NAND2X1 g34516(.A (u5_mem_b1_b_63 ), .B (n_7870), .Y (n_7912));
NAND2X1 g34517(.A (u5_mem_b1_b_64 ), .B (n_7870), .Y (n_7911));
NAND2X1 g34514(.A (u5_mem_b1_b_90 ), .B (n_7870), .Y (n_7914));
NAND2X1 g34515(.A (u5_mem_b1_b_62 ), .B (n_7870), .Y (n_7913));
NAND2X1 g39828(.A (u5_mem_b2_b_47 ), .B (n_12823), .Y (n_2243));
NAND2X1 g34636(.A (u6_mem_b2_b_40 ), .B (n_7758), .Y (n_7789));
NAND2X1 g36787(.A (n_1568), .B (n_1763), .Y (n_4064));
NAND2X1 g39704(.A (u4_mem_b1_b_79 ), .B (n_12265), .Y (n_4140));
NAND4X1 g36831(.A (n_11650), .B (n_11651), .C (n_2906), .D (n_11472),.Y (n_6777));
NOR2X1 g45677(.A (n_11672), .B (dma_ack_i_b6_b), .Y (n_12374));
NAND2X1 g45676(.A (dma_req_o_b6_b), .B (n_12370), .Y (n_12372));
NAND2X1 g39824(.A (u3_mem_b1_b_86 ), .B (n_3316), .Y (n_2938));
NOR2X1 g39707(.A (n_3117), .B (n_2702), .Y (n_3006));
INVX1 g42540(.A (u9_mem_b1_b ), .Y (n_6956));
INVX1 g36837(.A (n_6209), .Y (n_5726));
OAI21X1 g45675(.A0 (n_12371), .A1 (n_11672), .B0 (n_12372), .Y(n_12373));
NAND2X1 g39827(.A (n_11798), .B (u8_mem_b0_b_117 ), .Y (n_2935));
INVX2 g42860(.A (n_12634), .Y (n_6118));
INVX4 g45674(.A (n_12365), .Y (n_12369));
NOR2X1 g40038(.A (n_2772), .B (n_2182), .Y (n_2183));
NOR2X1 g39826(.A (n_3089), .B (n_2801), .Y (n_2937));
NOR2X1 g40036(.A (n_2470), .B (n_2829), .Y (n_1792));
NOR2X1 g40037(.A (n_2736), .B (n_2720), .Y (n_2809));
NOR2X1 g40034(.A (n_2470), .B (n_2707), .Y (n_2184));
NOR2X1 g40035(.A (n_2761), .B (n_2804), .Y (n_2811));
NOR2X1 g40032(.A (n_2043), .B (n_2741), .Y (n_2185));
NOR2X1 g40033(.A (n_2836), .B (n_2681), .Y (n_2812));
NOR2X1 g40030(.A (n_2742), .B (n_2735), .Y (n_2813));
NOR2X1 g40031(.A (n_2144), .B (n_2792), .Y (n_2186));
NAND2X1 g37159(.A (n_3910), .B (n_2241), .Y (n_6596));
NAND2X1 g37158(.A (n_3913), .B (n_2357), .Y (n_6599));
NAND2X1 g37153(.A (n_3905), .B (n_2279), .Y (n_6473));
NAND2X1 g37152(.A (n_2633), .B (n_4239), .Y (n_6646));
NAND2X1 g37151(.A (n_4618), .B (n_3195), .Y (n_6891));
NAND2X1 g37150(.A (n_4613), .B (n_2255), .Y (n_6906));
NAND2X1 g37157(.A (n_3920), .B (n_2280), .Y (n_6602));
NAND2X1 g37156(.A (n_2521), .B (n_2236), .Y (n_5997));
NAND2X1 g37155(.A (n_4615), .B (n_3347), .Y (n_6899));
NAND2X1 g37154(.A (n_2552), .B (n_2303), .Y (n_6017));
OAI21X1 g33466(.A0 (n_4513), .A1 (n_8393), .B0 (n_8109), .Y (n_8394));
XOR2X1 g36202(.A (n_4088), .B (n_1282), .Y (n_4089));
INVX2 g45672(.A (n_12364), .Y (n_12365));
NOR2X1 g39820(.A (n_3486), .B (n_2707), .Y (n_2941));
INVX1 g45671(.A (n_12365), .Y (n_12366));
INVX4 g40726(.A (n_940), .Y (n_2364));
NOR2X1 g39823(.A (n_4996), .B (n_2741), .Y (n_2939));
MX2X1 g33090(.A (n_56), .B (wb_din_670), .S0 (n_8643), .Y (n_8654));
NAND2X1 g39822(.A (in_slt_403), .B (n_3415), .Y (n_2940));
INVX8 g41259(.A (n_914), .Y (n_6649));
INVX1 g41255(.A (n_840), .Y (n_1142));
CLKBUFX1 g41254(.A (n_1142), .Y (n_4616));
MX2X1 g33099(.A (n_71), .B (wb_din_663), .S0 (n_8643), .Y (n_8641));
CLKBUFX3 g41253(.A (n_840), .Y (n_1143));
INVX8 g41252(.A (n_1143), .Y (n_2368));
OAI21X1 g31007(.A0 (n_5364), .A1 (n_10450), .B0 (n_10009), .Y(n_10694));
OAI21X1 g31006(.A0 (n_5521), .A1 (n_10679), .B0 (n_10011), .Y(n_10695));
OAI21X1 g31005(.A0 (n_5576), .A1 (n_10450), .B0 (n_10012), .Y(n_10697));
OAI21X1 g31004(.A0 (n_5578), .A1 (n_10450), .B0 (n_10013), .Y(n_10699));
OAI21X1 g31003(.A0 (n_5351), .A1 (n_10738), .B0 (n_10014), .Y(n_10700));
OAI21X1 g31002(.A0 (n_5366), .A1 (n_10747), .B0 (n_10015), .Y(n_10701));
OAI21X1 g31001(.A0 (n_5346), .A1 (n_10738), .B0 (n_10016), .Y(n_10702));
OAI21X1 g31000(.A0 (n_5348), .A1 (n_10738), .B0 (n_10017), .Y(n_10703));
NAND2X1 g39908(.A (n_3339), .B (in_slt_426), .Y (n_5292));
INVX1 g42780(.A (u11_mem_b2_b_110 ), .Y (n_277));
INVX1 g42786(.A (u11_mem_b1_b_121 ), .Y (n_6492));
OAI21X1 g31009(.A0 (n_5517), .A1 (n_10679), .B0 (n_10007), .Y(n_10691));
OAI21X1 g31008(.A0 (n_5519), .A1 (n_10450), .B0 (n_10008), .Y(n_10693));
CLKBUFX2 g45561(.A (n_12167), .Y (n_12168));
INVX4 g45560(.A (n_12168), .Y (n_12169));
XOR2X1 g40402(.A (n_1424), .B (n_1924), .Y (n_5620));
INVX1 g41784(.A (n_12332), .Y (n_754));
INVX1 g35041(.A (n_7414), .Y (n_9326));
INVX1 g41781(.A (n_754), .Y (n_907));
NAND2X1 g39909(.A (n_11798), .B (u8_mem_b0_b_103 ), .Y (n_11455));
INVX1 g41789(.A (u11_mem_b3_b_82 ), .Y (n_5500));
INVX1 g41788(.A (u11_mem_b1_b_136 ), .Y (n_1650));
INVX1 g41078(.A (n_818), .Y (n_819));
INVX4 g33351(.A (n_10483), .Y (n_10583));
OR2X1 g29972(.A (u13_ints_r_b2_b ), .B (oc0_int_set), .Y (n_10831));
INVX4 g41073(.A (n_1214), .Y (n_1575));
INVX8 g33355(.A (n_9873), .Y (n_10483));
NAND2X1 g41077(.A (n_3559), .B (n_771), .Y (n_923));
NAND2X2 g41076(.A (u11_rp_b1_b ), .B (n_487), .Y (n_1214));
MX2X1 g31263(.A (n_5479), .B (n_1704), .S0 (n_10303), .Y (n_10157));
MX2X1 g31262(.A (n_5481), .B (n_1701), .S0 (n_10303), .Y (n_10158));
MX2X1 g31261(.A (n_5482), .B (n_1733), .S0 (n_10308), .Y (n_10159));
MX2X1 g31260(.A (n_5483), .B (n_1562), .S0 (n_10308), .Y (n_10160));
MX2X1 g31267(.A (n_6860), .B (n_6859), .S0 (n_10267), .Y (n_10152));
OR2X1 g29970(.A (u13_ints_r_b14_b ), .B (oc4_int_set), .Y (n_10833));
MX2X1 g31265(.A (n_5475), .B (n_1724), .S0 (n_10308), .Y (n_10155));
MX2X1 g31264(.A (n_5477), .B (n_1728), .S0 (n_10308), .Y (n_10156));
NOR2X1 g39992(.A (n_2218), .B (n_2744), .Y (n_2212));
MX2X1 g31269(.A (n_5487), .B (n_1716), .S0 (n_10267), .Y (n_10150));
MX2X1 g31268(.A (n_5473), .B (n_2507), .S0 (n_10267), .Y (n_10151));
AOI21X1 g38031(.A0 (u3_mem_b3_b_149 ), .A1 (n_5138), .B0 (n_3358), .Y(n_5142));
AOI21X1 g35479(.A0 (i4_dout_611), .A1 (n_7468), .B0 (n_7140), .Y(n_7330));
OR2X1 g41631(.A (n_11777), .B (n_518), .Y (n_807));
XOR2X1 g40400(.A (n_1417), .B (n_11585), .Y (n_5618));
NOR2X1 g39888(.A (n_3089), .B (n_2720), .Y (n_2902));
NOR2X1 g35652(.A (u11_rp_b0_b ), .B (i6_re), .Y (n_6709));
NOR2X1 g40979(.A (n_1921), .B (n_1421), .Y (n_1422));
NAND3X1 g30112(.A (n_10985), .B (n_9996), .C (n_10331), .Y (n_10986));
INVX1 g41630(.A (n_807), .Y (n_1230));
MX2X1 g40433(.A (crac_din_705), .B (in_slt_844), .S0 (n_1036), .Y(n_1030));
AOI21X1 g38458(.A0 (u3_mem_b2_b_41 ), .A1 (n_4519), .B0 (n_2097), .Y(n_4325));
AOI22X1 g40407(.A0 (u13_intm_r_b10_b ), .A1 (u13_ints_r_b10_b ), .B0(u13_intm_r_b9_b ), .B1 (u13_ints_r_b9_b ), .Y (n_574));
OR2X1 g30110(.A (u13_ints_r_b23_b ), .B (ic1_int_set), .Y (n_9692));
NAND2X1 g39887(.A (n_12826), .B (u3_mem_b0_b_118 ), .Y (n_2903));
NOR2X1 g39904(.A (n_3453), .B (n_2801), .Y (n_2890));
AOI21X1 g35471(.A0 (i4_dout_615), .A1 (n_7468), .B0 (n_7136), .Y(n_7333));
OAI21X1 g31786(.A0 (n_5447), .A1 (n_9564), .B0 (n_9752), .Y (n_9964));
NOR2X1 g35476(.A (i4_empty), .B (i4_re), .Y (n_7148));
OAI21X1 g31039(.A0 (n_5318), .A1 (n_10820), .B0 (n_10370), .Y(n_10873));
INVX2 g40721(.A (n_941), .Y (n_1176));
NOR2X1 g35477(.A (i6_empty), .B (i6_re), .Y (n_7018));
OAI21X1 g31036(.A0 (n_5412), .A1 (n_10820), .B0 (n_10373), .Y(n_10877));
MX2X1 g40434(.A (crac_din_706), .B (in_slt_845), .S0 (n_1036), .Y(n_1083));
OAI21X1 g31789(.A0 (crac_out_876), .A1 (n_8486), .B0 (n_9794), .Y(n_10339));
NAND3X1 g40406(.A (n_594), .B (wb_addr_i_b3_b), .C (wb_addr_i_b4_b), .Y(n_1231));
MX2X1 g40428(.A (crac_din_699), .B (in_slt_838), .S0 (n_1036), .Y(n_1037));
NAND2X1 g39886(.A (u5_mem_b1_b_69 ), .B (n_3236), .Y (n_12030));
INVX1 g42297(.A (u9_mem_b0_b_180 ), .Y (n_1716));
INVX1 g42254(.A (u3_wp_b2_b ), .Y (n_214));
INVX1 g42250(.A (u10_mem_b2_b_118 ), .Y (n_1863));
INVX1 g42520(.A (u9_mem_b0_b_162 ), .Y (n_6392));
INVX1 g42521(.A (u10_mem_b2_b_106 ), .Y (n_256));
INVX1 g40405(.A (n_1231), .Y (n_2575));
NOR2X1 g39885(.A (n_3089), .B (n_2818), .Y (n_2905));
INVX1 g42528(.A (u10_mem_b1_b_136 ), .Y (n_313));
INVX2 g43124(.A (u4_rp_b0_b ), .Y (n_6824));
OAI21X1 g45806(.A0 (n_5720), .A1 (n_6995), .B0 (n_5860), .Y(n_12521));
INVX1 g43129(.A (u9_mem_b1_b_147 ), .Y (n_206));
INVX2 g43128(.A (u4_rp_b0_b ), .Y (n_145));
NAND2X1 g45803(.A (n_5869), .B (n_3559), .Y (n_12517));
AOI21X1 g35588(.A0 (n_6320), .A1 (n_5776), .B0 (n_7267), .Y (n_7269));
AOI21X1 g35589(.A0 (n_6319), .A1 (n_5775), .B0 (n_7267), .Y (n_7268));
NOR2X1 g35586(.A (n_1206), .B (i4_re), .Y (n_6712));
NOR2X1 g35587(.A (n_1039), .B (i4_re), .Y (n_6711));
AOI21X1 g35585(.A0 (n_6321), .A1 (n_6132), .B0 (n_7324), .Y (n_7270));
NOR2X1 g39003(.A (n_2732), .B (n_1488), .Y (n_1504));
AOI21X1 g35583(.A0 (n_6304), .A1 (n_5757), .B0 (n_7214), .Y (n_7271));
AOI21X1 g35580(.A0 (n_11541), .A1 (n_11542), .B0 (n_12145), .Y(n_7319));
AOI21X1 g35581(.A0 (n_6323), .A1 (n_6125), .B0 (n_12145), .Y(n_7273));
NAND2X1 g36859(.A (n_1691), .B (n_3927), .Y (n_5391));
NOR2X1 g36858(.A (n_5422), .B (n_6594), .Y (n_4819));
NAND2X1 g36855(.A (n_2504), .B (n_1692), .Y (n_4342));
NAND4X1 g36854(.A (n_11666), .B (n_11667), .C (n_3376), .D (n_2634),.Y (n_6254));
NAND2X1 g36857(.A (n_4078), .B (n_1249), .Y (n_5392));
NOR2X1 g36856(.A (n_5418), .B (n_6594), .Y (n_4820));
INVX1 g36851(.A (n_12530), .Y (n_5725));
NAND4X1 g36850(.A (n_4208), .B (n_3388), .C (n_2304), .D (n_4256), .Y(n_6800));
INVX1 g36853(.A (n_6254), .Y (n_5724));
INVX4 g34989(.A (n_7423), .Y (n_8101));
NAND2X1 g39883(.A (u4_mem_b2_b_42 ), .B (n_12091), .Y (n_2906));
NAND2X1 g39900(.A (u8_mem_b2_b_37 ), .B (n_2366), .Y (n_11450));
INVX2 g34983(.A (n_7423), .Y (n_8097));
AOI22X1 g37625(.A0 (n_6935), .A1 (n_1835), .B0 (n_6951), .B1(n_1760), .Y (n_1751));
NOR2X1 g39882(.A (n_2786), .B (n_1488), .Y (n_1322));
AOI22X1 g37624(.A0 (n_2502), .A1 (n_6864), .B0 (n_6954), .B1(n_1859), .Y (n_1752));
AOI22X1 g37627(.A0 (n_2502), .A1 (n_174), .B0 (n_1748), .B1 (n_1859),.Y (n_1749));
AOI22X1 g37626(.A0 (n_204), .A1 (n_1859), .B0 (n_6089), .B1 (n_1760),.Y (n_1750));
INVX1 g41001(.A (n_1416), .Y (n_2832));
AOI22X1 g37621(.A0 (n_6635), .A1 (n_1835), .B0 (n_6581), .B1(n_1760), .Y (n_1758));
NAND4X1 g33322(.A (n_6047), .B (n_2645), .C (n_7496), .D (n_968), .Y(n_9451));
AOI22X1 g37620(.A0 (n_2502), .A1 (n_6396), .B0 (n_6528), .B1(n_1859), .Y (n_1759));
AOI22X1 g40409(.A0 (u13_intm_r_b7_b ), .A1 (u13_ints_r_b7_b ), .B0(u13_intm_r_b8_b ), .B1 (u13_ints_r_b8_b ), .Y (n_543));
NOR2X1 g39881(.A (n_3453), .B (n_2794), .Y (n_2907));
INVX1 g41003(.A (n_1416), .Y (n_2742));
AOI22X1 g37623(.A0 (n_2502), .A1 (n_6866), .B0 (n_6922), .B1(n_1760), .Y (n_1753));
AOI22X1 g37622(.A0 (n_1756), .A1 (n_1755), .B0 (n_1754), .B1(n_1643), .Y (n_1757));
INVX1 g41005(.A (n_1416), .Y (n_2788));
INVX2 g41007(.A (n_1016), .Y (n_1416));
AOI22X1 g40408(.A0 (u13_intm_r_b2_b ), .A1 (u13_ints_r_b2_b ), .B0(u13_intm_r_b4_b ), .B1 (u13_ints_r_b4_b ), .Y (n_549));
NAND2X1 g39880(.A (u8_mem_b2_b_41 ), .B (n_2362), .Y (n_1867));
NAND2X2 g41008(.A (n_1424), .B (n_626), .Y (n_1016));
INVX2 g41009(.A (n_928), .Y (n_6259));
NAND2X1 g34239(.A (u3_mem_b1_b_89 ), .B (n_8101), .Y (n_8167));
NAND2X1 g34238(.A (u8_mem_b2_b_37 ), .B (n_7976), .Y (n_8168));
OAI21X1 g33517(.A0 (n_4462), .A1 (n_9346), .B0 (n_8042), .Y (n_8330));
OAI21X1 g33516(.A0 (n_4463), .A1 (n_9346), .B0 (n_8044), .Y (n_8332));
NAND2X1 g34235(.A (u3_mem_b1_b_88 ), .B (n_8101), .Y (n_8172));
NAND2X1 g34234(.A (u8_mem_b2_b_33 ), .B (n_7976), .Y (n_8173));
OAI21X1 g33513(.A0 (n_4465), .A1 (n_9349), .B0 (n_8048), .Y (n_8338));
OAI21X1 g33512(.A0 (n_4467), .A1 (n_8333), .B0 (n_8049), .Y (n_8340));
OAI21X1 g33511(.A0 (n_4469), .A1 (n_8333), .B0 (n_8051), .Y (n_8341));
OAI21X1 g33510(.A0 (n_4470), .A1 (n_9346), .B0 (n_8052), .Y (n_8342));
NOR2X1 g41303(.A (n_670), .B (n_921), .Y (n_690));
NAND2X2 g41302(.A (n_691), .B (n_12281), .Y (n_692));
AOI21X1 g35955(.A0 (n_6972), .A1 (oc1_cfg_976), .B0 (n_5795), .Y(n_6973));
INVX2 g37526(.A (n_1779), .Y (n_6686));
NAND3X1 g37527(.A (n_1132), .B (wb_addr_i_b6_b), .C (n_593), .Y(n_1779));
BUFX3 g40770(.A (n_945), .Y (n_4533));
NAND2X1 g37528(.A (n_5645), .B (n_2968), .Y (n_4653));
NOR2X1 g37529(.A (n_5309), .B (n_6649), .Y (n_4652));
OAI21X1 g33632(.A0 (n_5013), .A1 (n_9212), .B0 (n_7910), .Y (n_9278));
OAI21X1 g33633(.A0 (n_5012), .A1 (n_9307), .B0 (n_7909), .Y (n_9277));
OAI21X1 g33630(.A0 (n_5015), .A1 (n_9286), .B0 (n_7912), .Y (n_9281));
OAI21X1 g33631(.A0 (n_5014), .A1 (n_9286), .B0 (n_7911), .Y (n_9280));
OAI21X1 g33636(.A0 (n_4379), .A1 (n_9286), .B0 (n_7904), .Y (n_9274));
OAI21X1 g33637(.A0 (n_4377), .A1 (n_9288), .B0 (n_7903), .Y (n_9273));
OAI21X1 g33634(.A0 (n_5141), .A1 (n_9286), .B0 (n_7908), .Y (n_9276));
OAI21X1 g33826(.A0 (n_4895), .A1 (n_9036), .B0 (n_7698), .Y (n_9040));
INVX1 g40775(.A (n_1172), .Y (n_2120));
OAI21X1 g33638(.A0 (n_4376), .A1 (n_9307), .B0 (n_7902), .Y (n_9272));
OAI21X1 g33639(.A0 (n_4375), .A1 (n_9307), .B0 (n_7901), .Y (n_9270));
OAI21X1 g33825(.A0 (n_4911), .A1 (n_9010), .B0 (n_7699), .Y (n_9041));
OAI21X1 g35950(.A0 (n_5528), .A1 (n_6981), .B0 (n_5799), .Y (n_6976));
NAND2X1 g38981(.A (u8_mem_b3_b_125 ), .B (n_2468), .Y (n_2382));
OAI21X1 g33824(.A0 (n_4896), .A1 (n_9038), .B0 (n_7701), .Y (n_9042));
NAND2X1 g39218(.A (n_11798), .B (u8_mem_b0_b_120 ), .Y (n_3360));
NAND2X1 g38980(.A (u8_mem_b3_b_146 ), .B (n_2468), .Y (n_2383));
NAND2X1 g34291(.A (u3_mem_b2_b_35 ), .B (n_8101), .Y (n_8107));
INVX1 g42798(.A (u11_mem_b2_b_94 ), .Y (n_6530));
NAND2X1 g39219(.A (n_12747), .B (u4_rp_b3_b ), .Y (n_5466));
NAND2X1 g38983(.A (u8_mem_b3_b_141 ), .B (n_2468), .Y (n_2380));
OAI21X1 g33822(.A0 (n_4897), .A1 (n_9043), .B0 (n_7703), .Y (n_9045));
INVX1 g40779(.A (n_1172), .Y (n_2083));
NAND2X1 g38982(.A (u8_mem_b3_b_126 ), .B (n_2468), .Y (n_2381));
OAI21X1 g33821(.A0 (n_4964), .A1 (n_9034), .B0 (n_7704), .Y (n_9046));
INVX1 g40778(.A (n_1172), .Y (n_2071));
INVX1 g38985(.A (n_1132), .Y (n_1133));
OAI21X1 g33820(.A0 (n_4899), .A1 (n_9010), .B0 (n_7705), .Y (n_9047));
AOI21X1 g38530(.A0 (u7_mem_b3_b_134 ), .A1 (n_5145), .B0 (n_3342), .Y(n_4874));
AOI21X1 g38531(.A0 (u3_mem_b2_b_44 ), .A1 (n_4519), .B0 (n_1934), .Y(n_4296));
AOI21X1 g38532(.A0 (u4_mem_b1_b_68 ), .A1 (n_4507), .B0 (n_2107), .Y(n_4295));
AOI21X1 g38533(.A0 (u7_mem_b2_b_36 ), .A1 (n_4509), .B0 (n_2181), .Y(n_4294));
AOI21X1 g38534(.A0 (u3_mem_b2_b_32 ), .A1 (n_4533), .B0 (n_1950), .Y(n_4293));
AOI21X1 g38535(.A0 (u3_mem_b3_b_131 ), .A1 (n_5133), .B0 (n_3090), .Y(n_4873));
AOI21X1 g38536(.A0 (u7_mem_b2_b_35 ), .A1 (n_4540), .B0 (n_1942), .Y(n_4292));
AOI21X1 g38537(.A0 (u3_mem_b1_b_80 ), .A1 (n_5148), .B0 (n_2695), .Y(n_4872));
AOI21X1 g38538(.A0 (u3_mem_b3_b_132 ), .A1 (n_5138), .B0 (n_2858), .Y(n_4871));
AOI21X1 g38539(.A0 (u8_mem_b3_b_138 ), .A1 (n_3879), .B0 (n_1457), .Y(n_3843));
AOI21X1 g38234(.A0 (u4_mem_b3_b_130 ), .A1 (n_5102), .B0 (n_3007), .Y(n_5064));
NOR2X1 g39213(.A (n_3453), .B (n_2782), .Y (n_3364));
MX2X1 g33184(.A (wb_din_669), .B (oc5_cfg_1014), .S0 (n_8202), .Y(n_8184));
MX2X1 g33180(.A (wb_din_665), .B (n_8188), .S0 (n_8202), .Y (n_8189));
MX2X1 g33181(.A (wb_din_666), .B (n_4701), .S0 (n_8202), .Y (n_8187));
MX2X1 g33182(.A (wb_din_667), .B (oc4_cfg_1010), .S0 (n_8202), .Y(n_8186));
MX2X1 g33183(.A (wb_din_668), .B (n_8182), .S0 (n_8202), .Y (n_8185));
AOI21X1 g38238(.A0 (u6_mem_b3_b_151 ), .A1 (n_5100), .B0 (n_2998), .Y(n_5062));
INVX4 g40522(.A (wb_din_681), .Y (n_2729));
NOR2X1 g39645(.A (n_2804), .B (n_1488), .Y (n_1478));
AOI21X1 g37995(.A0 (u6_mem_b2_b_55 ), .A1 (n_4544), .B0 (n_2082), .Y(n_4545));
NAND2X1 g36693(.A (n_5539), .B (n_6118), .Y (n_6095));
OAI21X1 g36691(.A0 (n_5455), .A1 (n_5456), .B0 (n_6118), .Y (n_6097));
OAI21X1 g36690(.A0 (n_5451), .A1 (n_5457), .B0 (n_6118), .Y (n_6099));
OAI21X1 g36697(.A0 (n_5194), .A1 (n_5193), .B0 (n_634), .Y (n_5757));
NAND2X1 g36694(.A (n_5699), .B (n_6118), .Y (n_6761));
OAI21X1 g36698(.A0 (n_4627), .A1 (n_5191), .B0 (n_634), .Y (n_5756));
NAND2X1 g39644(.A (u6_mem_b1_b_80 ), .B (n_4253), .Y (n_4154));
NAND2X1 g45782(.A (n_12411), .B (n_6118), .Y (n_12496));
NAND2X1 g45781(.A (n_12634), .B (n_6228), .Y (n_12495));
AOI21X1 g45780(.A0 (n_12495), .A1 (n_12496), .B0 (n_12640), .Y(n_12499));
CLKBUFX3 g45787(.A (n_12502), .Y (n_12503));
CLKBUFX3 g45786(.A (n_12503), .Y (n_12504));
OAI21X1 g45785(.A0 (n_5542), .A1 (n_7088), .B0 (n_5819), .Y(n_12500));
OR2X1 g45789(.A (n_11528), .B (n_8663), .Y (n_12501));
INVX1 g45788(.A (n_12501), .Y (n_12502));
NOR2X1 g30725(.A (n_10810), .B (n_11144), .Y (n_11112));
OAI21X1 g30724(.A0 (n_5436), .A1 (n_9651), .B0 (n_9650), .Y (n_9652));
NOR2X1 g30727(.A (n_10657), .B (n_11126), .Y (n_11004));
NOR2X1 g30726(.A (n_10773), .B (n_11126), .Y (n_11005));
NOR2X1 g30721(.A (n_10774), .B (n_11131), .Y (n_11007));
NOR2X1 g30720(.A (n_10811), .B (n_11086), .Y (n_11113));
NOR2X1 g30722(.A (n_10659), .B (n_11131), .Y (n_11006));
OR2X1 g30729(.A (n_10404), .B (n_11136), .Y (n_11002));
OR2X1 g30728(.A (n_10405), .B (n_12589), .Y (n_11512));
BUFX3 g35009(.A (o3_we), .Y (n_7423));
INVX2 g35002(.A (n_7423), .Y (n_8856));
CLKBUFX1 g35000(.A (o3_we), .Y (n_7424));
NAND2X1 g39691(.A (u6_mem_b1_b_79 ), .B (n_12169), .Y (n_4143));
MX2X1 g36079(.A (n_6507), .B (n_6465), .S0 (n_995), .Y (n_6508));
MX2X1 g36078(.A (n_5994), .B (n_5993), .S0 (n_5312), .Y (n_5995));
MX2X1 g36077(.A (n_6511), .B (n_6510), .S0 (n_995), .Y (n_6512));
MX2X1 g36076(.A (n_6515), .B (n_6514), .S0 (n_6502), .Y (n_6516));
MX2X1 g36075(.A (n_6517), .B (n_6473), .S0 (n_6502), .Y (n_6518));
MX2X1 g36074(.A (n_6519), .B (n_6478), .S0 (n_6502), .Y (n_6520));
MX2X1 g36073(.A (n_6522), .B (n_6521), .S0 (n_6502), .Y (n_6523));
MX2X1 g36072(.A (n_6497), .B (n_6524), .S0 (n_6649), .Y (n_6525));
MX2X1 g36071(.A (n_6526), .B (n_6579), .S0 (n_6475), .Y (n_6527));
MX2X1 g36070(.A (n_6873), .B (n_6883), .S0 (n_6898), .Y (n_6874));
NAND2X1 g37449(.A (u13_ints_r_b11_b ), .B (n_3979), .Y (n_3980));
INVX1 g42068(.A (u11_mem_b3_b_68 ), .Y (n_6604));
AND2X1 g41355(.A (u11_wp_b0_b ), .B (u11_wp_b1_b ), .Y (n_512));
INVX1 g42062(.A (u8_wp_b0_b ), .Y (n_58));
INVX1 g42060(.A (u9_mem_b1_b_149 ), .Y (n_1715));
INVX1 g42067(.A (oc1_int_set_709), .Y (n_540));
INVX1 g42065(.A (u11_mem_b0_b_166 ), .Y (n_5951));
NAND2X1 g39641(.A (n_12369), .B (u6_mem_b0_b_110 ), .Y (n_3041));
NAND3X1 g34712(.A (n_5588), .B (n_5788), .C (n_863), .Y (n_1885));
NAND2X1 g39698(.A (u4_mem_b2_b_50 ), .B (n_12091), .Y (n_3013));
OAI21X1 g35919(.A0 (n_5693), .A1 (n_7080), .B0 (n_6197), .Y (n_7079));
OAI21X1 g35911(.A0 (n_5726), .A1 (n_7088), .B0 (n_6774), .Y (n_7182));
OAI21X1 g35910(.A0 (n_5690), .A1 (n_7088), .B0 (n_6208), .Y (n_7084));
OAI21X1 g35913(.A0 (n_6072), .A1 (n_7088), .B0 (n_6206), .Y (n_7179));
OAI21X1 g35912(.A0 (n_5688), .A1 (n_7088), .B0 (n_6772), .Y (n_7181));
OAI21X1 g35914(.A0 (n_6070), .A1 (n_7088), .B0 (n_6771), .Y (n_7178));
OAI21X1 g35917(.A0 (n_5696), .A1 (n_7080), .B0 (n_6199), .Y (n_7081));
NAND2X1 g39640(.A (u8_mem_b1_b ), .B (n_12295), .Y (n_11468));
INVX1 g41826(.A (dma_req_o_b5_b), .Y (n_284));
NAND2X1 g39643(.A (u6_mem_b2_b_49 ), .B (n_3423), .Y (n_3038));
INVX1 g41827(.A (u9_mem_b2_b_107 ), .Y (n_1744));
NAND2X1 g34758(.A (u7_mem_b2_b_45 ), .B (n_7651), .Y (n_7676));
NAND2X1 g34759(.A (u7_mem_b2_b_46 ), .B (n_7651), .Y (n_7675));
BUFX3 g40900(.A (n_2553), .Y (n_2544));
NAND2X1 g34750(.A (u7_mem_b2_b ), .B (n_7651), .Y (n_7684));
NAND2X1 g34751(.A (u7_mem_b2_b_38 ), .B (n_7651), .Y (n_7683));
NAND2X1 g34752(.A (u7_mem_b2_b_39 ), .B (n_7651), .Y (n_7682));
NAND2X1 g34753(.A (u7_mem_b2_b_40 ), .B (n_7651), .Y (n_7681));
NAND2X1 g34754(.A (u7_mem_b2_b_41 ), .B (n_7651), .Y (n_7680));
NAND2X1 g34755(.A (u7_mem_b2_b_42 ), .B (n_7651), .Y (n_7679));
NAND2X1 g34756(.A (u7_mem_b2_b_43 ), .B (n_7651), .Y (n_7678));
NAND2X1 g34757(.A (u7_mem_b2_b_44 ), .B (n_7651), .Y (n_7677));
AND2X1 g35322(.A (n_1136), .B (n_6718), .Y (n_11887));
NOR2X1 g39252(.A (n_3486), .B (n_2716), .Y (n_3343));
NAND2X1 g39253(.A (u5_mem_b2_b_37 ), .B (n_12823), .Y (n_2337));
NAND2X1 g39250(.A (u8_mem_b2_b_36 ), .B (n_2362), .Y (n_2338));
NAND2X1 g39251(.A (u3_mem_b1_b_62 ), .B (n_3316), .Y (n_3701));
INVX1 g39256(.A (n_5309), .Y (n_4207));
NAND2X1 g39257(.A (n_4560), .B (in_slt_454), .Y (n_5309));
NOR2X1 g39255(.A (n_4961), .B (n_2681), .Y (n_3342));
NAND2X1 g39258(.A (u3_mem_b2_b_39 ), .B (n_12619), .Y (n_3341));
NAND2X1 g39259(.A (n_2325), .B (in_slt_442), .Y (n_2472));
NAND2X1 g34534(.A (u5_mem_b2_b_29 ), .B (n_7870), .Y (n_7893));
NAND2X1 g34535(.A (u5_mem_b2_b_48 ), .B (n_7870), .Y (n_7892));
NAND2X1 g34536(.A (u5_mem_b2_b_49 ), .B (n_7870), .Y (n_7891));
NAND2X1 g34537(.A (u5_mem_b2_b_50 ), .B (n_7870), .Y (n_7890));
NAND2X1 g34530(.A (u5_mem_b2_b_44 ), .B (n_7870), .Y (n_7897));
NAND2X1 g34531(.A (u5_mem_b2_b_45 ), .B (n_7870), .Y (n_7896));
NAND2X1 g34532(.A (u5_mem_b2_b_46 ), .B (n_7870), .Y (n_7895));
NAND2X1 g34533(.A (u5_mem_b2_b_47 ), .B (n_7870), .Y (n_7894));
AND2X1 g35323(.A (n_1105), .B (n_6720), .Y (n_11888));
INVX1 g41868(.A (u9_mem_b0_b_156 ), .Y (n_6847));
NAND2X1 g34538(.A (u5_mem_b2_b_51 ), .B (n_7870), .Y (n_7889));
NAND2X1 g34539(.A (u5_mem_b2_b_52 ), .B (n_7870), .Y (n_7888));
NAND2X1 g34618(.A (u6_mem_b1_b_86 ), .B (n_7758), .Y (n_7807));
NAND2X1 g39646(.A (n_12204), .B (u6_mem_b0_b_111 ), .Y (n_3037));
NOR2X1 g40045(.A (n_2759), .B (n_3008), .Y (n_2806));
NOR2X1 g39999(.A (n_2736), .B (n_2767), .Y (n_2826));
NAND2X1 g39727(.A (u6_mem_b2_b_30 ), .B (n_2285), .Y (n_11515));
NAND2X1 g34797(.A (u7_mem_b3_b_145 ), .B (n_7651), .Y (n_7636));
NAND2X1 g39648(.A (n_3339), .B (in_slt_435), .Y (n_5284));
NOR2X1 g41614(.A (u3_rp_b3_b ), .B (u3_wp_b2_b ), .Y (n_477));
NAND2X1 g39723(.A (n_4560), .B (in_slt_452), .Y (n_5321));
OAI21X1 g33441(.A0 (n_3864), .A1 (n_8453), .B0 (n_8137), .Y (n_8422));
NOR2X1 g40018(.A (n_2749), .B (n_2790), .Y (n_2817));
NAND2X1 g40019(.A (n_4502), .B (n_4499), .Y (n_1454));
NOR2X1 g40010(.A (n_2696), .B (n_2818), .Y (n_2821));
NOR2X1 g40011(.A (n_2735), .B (n_2067), .Y (n_2202));
NOR2X1 g40012(.A (n_2818), .B (n_1985), .Y (n_2201));
NOR2X1 g40013(.A (n_2216), .B (n_2792), .Y (n_2199));
AOI21X1 g40014(.A0 (oc1_cfg_974), .A1 (in_slt_752), .B0(u14_u1_full_empty_r), .Y (n_620));
NOR2X1 g40015(.A (n_2736), .B (n_2831), .Y (n_2820));
NOR2X1 g40016(.A (n_867), .B (n_2741), .Y (n_2198));
INVX4 g41611(.A (n_745), .Y (n_5102));
AOI22X1 g37332(.A0 (n_5277), .A1 (crac_out_867), .B0 (n_6972), .B1(n_3987), .Y (n_3989));
INVX4 g41610(.A (n_5102), .Y (n_1475));
NAND2X1 g39583(.A (n_12825), .B (u3_mem_b0_b_110 ), .Y (n_3082));
NOR2X1 g41613(.A (u13_ints_r_b19_b ), .B (n_525), .Y (n_580));
NOR2X1 g40858(.A (n_6821), .B (u6_rp_b3_b ), .Y (n_709));
INVX1 g40836(.A (n_1167), .Y (n_2054));
NOR2X1 g41612(.A (n_744), .B (n_444), .Y (n_745));
INVX2 g41271(.A (n_841), .Y (n_1055));
AOI22X1 g37842(.A0 (n_1756), .A1 (n_6355), .B0 (n_6492), .B1(n_1643), .Y (n_1579));
INVX1 g40837(.A (n_1167), .Y (n_2133));
OAI21X1 g31061(.A0 (n_5285), .A1 (n_10450), .B0 (n_9977), .Y(n_10668));
OAI21X1 g31060(.A0 (n_4792), .A1 (n_10679), .B0 (n_9978), .Y(n_10666));
OAI21X1 g31063(.A0 (n_5583), .A1 (n_10880), .B0 (n_10357), .Y(n_10857));
OAI21X1 g31062(.A0 (n_5581), .A1 (n_10880), .B0 (n_10358), .Y(n_10858));
OAI21X1 g31065(.A0 (n_5362), .A1 (n_10450), .B0 (n_9976), .Y(n_10664));
OAI21X1 g31064(.A0 (n_5495), .A1 (n_10880), .B0 (n_10356), .Y(n_10856));
OAI21X1 g31067(.A0 (n_5489), .A1 (n_10820), .B0 (n_10354), .Y(n_10854));
OAI21X1 g31066(.A0 (n_5527), .A1 (n_10820), .B0 (n_10355), .Y(n_10855));
OAI21X1 g31069(.A0 (n_5491), .A1 (n_10880), .B0 (n_10353), .Y(n_10853));
OAI21X1 g31068(.A0 (n_5349), .A1 (n_10450), .B0 (n_9975), .Y(n_10665));
INVX4 g40908(.A (n_1000), .Y (n_1643));
NAND2X1 g40909(.A (n_5), .B (u11_rp_b0_b ), .Y (n_1000));
NAND3X1 g33372(.A (n_1481), .B (n_6841), .C (n_7651), .Y (n_8175));
AND2X1 g33370(.A (n_9352), .B (u14_u6_en_out_l2), .Y (n_9447));
NAND2X1 g41055(.A (n_12581), .B (u5_rp_b1_b ), .Y (n_587));
INVX2 g41054(.A (n_587), .Y (n_1035));
INVX1 g33379(.A (n_9564), .Y (n_9620));
INVX4 g41058(.A (n_1153), .Y (n_4097));
MX2X1 g33170(.A (wb_din_670), .B (oc5_cfg_1015), .S0 (n_8202), .Y(n_8203));
MX2X1 g31289(.A (n_6391), .B (n_6390), .S0 (n_10315), .Y (n_10133));
MX2X1 g31288(.A (n_6371), .B (n_6370), .S0 (n_10820), .Y (n_10818));
MX2X1 g31285(.A (n_6378), .B (n_6377), .S0 (n_10820), .Y (n_10821));
MX2X1 g31284(.A (n_6381), .B (n_6380), .S0 (n_10450), .Y (n_10449));
MX2X1 g31287(.A (n_6373), .B (n_6372), .S0 (n_10820), .Y (n_10819));
MX2X1 g31286(.A (n_6376), .B (n_6375), .S0 (n_10315), .Y (n_10134));
NAND2X1 g34543(.A (u5_mem_b2_b_56 ), .B (n_7870), .Y (n_7884));
MX2X1 g31280(.A (n_5960), .B (n_5959), .S0 (n_10137), .Y (n_10138));
MX2X1 g31283(.A (n_6383), .B (n_6382), .S0 (n_10450), .Y (n_10451));
MX2X1 g31282(.A (n_6385), .B (n_6384), .S0 (n_10137), .Y (n_10135));
AND2X1 g45469(.A (n_11659), .B (n_2233), .Y (n_11924));
INVX1 g45858(.A (u5_rp_b1_b ), .Y (n_12583));
INVX1 g45680(.A (dma_ack_i_b7_b), .Y (n_12375));
NAND2X1 g36486(.A (n_5859), .B (n_5876), .Y (n_5860));
NAND2X1 g36487(.A (n_5857), .B (n_5881), .Y (n_5858));
NAND2X1 g36484(.A (n_5869), .B (n_5876), .Y (n_5862));
NAND2X1 g36485(.A (n_5865), .B (n_5876), .Y (n_5861));
NAND2X1 g36482(.A (n_5863), .B (n_5876), .Y (n_5864));
NAND2X1 g36481(.A (n_5865), .B (n_1229), .Y (n_5866));
BUFX3 g40833(.A (n_867), .Y (n_4370));
INVX1 g42157(.A (u9_mem_b0_b_151 ), .Y (n_6859));
NAND2X1 g36488(.A (n_6239), .B (n_6141), .Y (n_6240));
NAND2X1 g36489(.A (n_3939), .B (n_4644), .Y (n_6756));
OAI21X1 g45462(.A0 (n_4631), .A1 (n_4630), .B0 (n_11912), .Y(n_11913));
NOR2X1 g41619(.A (n_1206), .B (n_5420), .Y (n_1207));
NAND2X1 g45460(.A (n_11911), .B (n_11913), .Y (n_11914));
INVX2 g41417(.A (n_737), .Y (n_1760));
NAND3X1 g45461(.A (n_6157), .B (n_6316), .C (n_12535), .Y (n_11911));
INVX1 g41828(.A (u10_mem_b2_b_99 ), .Y (n_6666));
NAND2X1 g45466(.A (n_11923), .B (n_11927), .Y (n_11928));
INVX2 g42156(.A (u3_rp_b1_b ), .Y (n_600));
INVX1 g41829(.A (u11_mem_b1_b_132 ), .Y (n_6507));
NAND2X1 g45467(.A (n_11925), .B (n_12357), .Y (n_11927));
NOR2X1 g30880(.A (n_10979), .B (n_5839), .Y (n_11135));
AOI21X1 g30881(.A0 (n_11617), .A1 (n_11618), .B0 (n_11036), .Y(n_11038));
NOR2X1 g30882(.A (n_10977), .B (n_5839), .Y (n_11134));
AOI21X1 g30883(.A0 (n_11619), .A1 (n_11620), .B0 (n_11036), .Y(n_11037));
AOI21X1 g30884(.A0 (n_12062), .A1 (n_12063), .B0 (n_5839), .Y(n_11035));
AOI21X1 g30885(.A0 (n_11627), .A1 (n_11628), .B0 (n_11033), .Y(n_11034));
AOI21X1 g30886(.A0 (n_11994), .A1 (n_11995), .B0 (n_5839), .Y(n_11032));
AOI21X1 g35619(.A0 (n_6782), .A1 (n_6305), .B0 (n_7256), .Y (n_7309));
AOI21X1 g30888(.A0 (n_11623), .A1 (n_11624), .B0 (n_11025), .Y(n_11029));
AOI21X1 g35617(.A0 (n_6766), .A1 (n_6307), .B0 (n_7256), .Y (n_7312));
AOI21X1 g35614(.A0 (n_5921), .A1 (n_6103), .B0 (n_7256), .Y (n_7249));
AOI21X1 g35612(.A0 (n_5922), .A1 (n_6139), .B0 (n_7256), .Y (n_7251));
AOI21X1 g35613(.A0 (n_5941), .A1 (n_6108), .B0 (n_7256), .Y (n_7250));
AOI21X1 g35610(.A0 (n_5923), .A1 (n_6138), .B0 (n_7256), .Y (n_7253));
AOI21X1 g35611(.A0 (n_6822), .A1 (n_6109), .B0 (n_7256), .Y (n_7314));
AOI21X1 g40404(.A0 (u9_rp_b2_b ), .A1 (u9_wp_b3_b ), .B0 (n_478), .Y(n_2621));
MX2X1 g36168(.A (n_5955), .B (n_6011), .S0 (n_6341), .Y (n_5956));
INVX1 g38773(.A (n_5442), .Y (n_1804));
INVX2 g42155(.A (n_600), .Y (n_656));
INVX1 g42502(.A (u9_mem_b1_b_132 ), .Y (n_6654));
MX2X1 g38771(.A (u7_mem_b0_b_108 ), .B (wb_din_678), .S0 (n_3622), .Y(n_3564));
INVX1 g42507(.A (n_1923), .Y (n_1012));
INVX1 g38776(.A (n_4851), .Y (n_3563));
NAND2X1 g39489(.A (n_12826), .B (u3_mem_b0_b ), .Y (n_12832));
ADDHX1 g38777(.A (u26_cnt_b0_b ), .B (u26_cnt_b1_b ), .CO (n_793), .S(n_794));
AOI21X1 g35559(.A0 (n_5585), .A1 (n_4721), .B0 (n_7353), .Y (n_7134));
ADDHX1 g38774(.A (u2_res_cnt_b1_b ), .B (u2_res_cnt_b0_b ), .CO(n_1277), .S (n_796));
INVX1 g42154(.A (n_656), .Y (n_1924));
AOI21X1 g35558(.A0 (n_5587), .A1 (n_4722), .B0 (n_7353), .Y (n_7135));
INVX1 g43107(.A (n_1203), .Y (n_605));
INVX1 g43103(.A (u11_mem_b1_b_134 ), .Y (n_5990));
INVX1 g43102(.A (u11_mem_b3_b_79 ), .Y (n_5490));
INVX1 g43100(.A (u10_mem_b1_b_145 ), .Y (n_143));
NAND2X1 g34426(.A (u4_mem_b2_b_34 ), .B (n_7984), .Y (n_7990));
NAND2X1 g36876(.A (n_1189), .B (n_2302), .Y (n_4036));
NAND4X1 g36875(.A (n_11465), .B (n_11466), .C (n_2509), .D (n_1881),.Y (n_5895));
INVX1 g36874(.A (n_5895), .Y (n_5567));
NAND4X1 g36873(.A (n_12038), .B (n_11503), .C (n_12039), .D (n_2453),.Y (n_6244));
NAND2X1 g36870(.A (n_3918), .B (n_1243), .Y (n_5385));
NAND2X1 g39063(.A (n_11798), .B (u8_mem_b0_b_96 ), .Y (n_11465));
NAND2X1 g39062(.A (u7_mem_b2_b_56 ), .B (n_12650), .Y (n_4234));
NAND2X1 g39065(.A (u6_mem_b2_b_55 ), .B (n_3423), .Y (n_3480));
NAND2X1 g39064(.A (u8_mem_b2_b_56 ), .B (n_2366), .Y (n_1915));
NAND2X1 g36879(.A (n_1678), .B (n_1675), .Y (n_4034));
NOR2X1 g36878(.A (n_2486), .B (n_2302), .Y (n_4035));
INVX1 g42152(.A (n_1924), .Y (n_1096));
NOR2X1 g39642(.A (n_3332), .B (n_2716), .Y (n_3040));
AOI21X1 g35555(.A0 (n_5590), .A1 (n_4686), .B0 (n_7353), .Y (n_7138));
AOI21X1 g35554(.A0 (n_5584), .A1 (n_4694), .B0 (n_7353), .Y (n_7139));
AOI21X1 g35556(.A0 (n_5789), .A1 (n_4727), .B0 (n_7353), .Y (n_7137));
NAND2X1 g34425(.A (u4_mem_b2_b_33 ), .B (n_7984), .Y (n_7991));
OAI21X1 g36639(.A0 (n_4607), .A1 (n_5219), .B0 (u4_rp_b0_b ), .Y(n_6125));
NAND2X1 g39807(.A (u7_mem_b1_b_60 ), .B (n_4130), .Y (n_4118));
INVX1 g42435(.A (n_8526), .Y (n_671));
NAND2X1 g34422(.A (u4_mem_b2_b_59 ), .B (n_7984), .Y (n_7994));
CLKBUFX1 g45356(.A (n_11578), .Y (n_11563));
NAND2X1 g39804(.A (u8_mem_b2_b ), .B (n_2362), .Y (n_2245));
INVX1 g43087(.A (in_slt_736), .Y (n_209));
NAND2X1 g34259(.A (u8_mem_b3_b_150 ), .B (n_7976), .Y (n_8143));
NAND2X1 g34258(.A (u3_mem_b2_b_38 ), .B (n_8141), .Y (n_8144));
NAND2X1 g34423(.A (u4_mem_b2_b_31 ), .B (n_7984), .Y (n_7993));
OAI21X1 g33571(.A0 (n_5114), .A1 (n_8318), .B0 (n_7986), .Y (n_8265));
NAND2X1 g34250(.A (u8_mem_b3_b_142 ), .B (n_7976), .Y (n_8152));
NAND2X1 g34253(.A (u8_mem_b3_b_145 ), .B (n_7976), .Y (n_8149));
OAI21X1 g33572(.A0 (n_5107), .A1 (n_8318), .B0 (n_7985), .Y (n_8264));
NAND2X1 g34255(.A (u8_mem_b3_b_147 ), .B (n_7976), .Y (n_8147));
NAND2X1 g34254(.A (u8_mem_b3_b_146 ), .B (n_7976), .Y (n_8148));
OAI21X1 g33577(.A0 (n_5098), .A1 (n_9349), .B0 (n_7978), .Y (n_9351));
NAND2X1 g34256(.A (u8_mem_b3_b_148 ), .B (n_7976), .Y (n_8146));
NAND2X1 g38919(.A (u3_mem_b3_b_129 ), .B (n_2463), .Y (n_2402));
AOI21X1 g38080(.A0 (u3_mem_b3_b_127 ), .A1 (n_5138), .B0 (n_3426), .Y(n_5121));
AOI21X1 g38081(.A0 (u8_mem_b3_b_145 ), .A1 (n_3879), .B0 (n_1496), .Y(n_3881));
AOI21X1 g38082(.A0 (u8_mem_b3_b_144 ), .A1 (n_3879), .B0 (n_1462), .Y(n_3880));
NAND2X1 g34420(.A (u4_mem_b2_b_30 ), .B (n_7984), .Y (n_7996));
NOR2X1 g37509(.A (n_5284), .B (n_6594), .Y (n_4658));
INVX1 g37058(.A (n_6150), .Y (n_5686));
NAND4X1 g37059(.A (n_12831), .B (n_12832), .C (n_2893), .D (n_1514),.Y (n_6150));
NOR2X1 g37504(.A (n_5355), .B (n_6594), .Y (n_4660));
NAND2X1 g37057(.A (n_2536), .B (n_1295), .Y (n_4806));
NAND4X1 g37054(.A (n_1516), .B (n_3523), .C (n_3483), .D (n_3553), .Y(n_5539));
NAND4X1 g37055(.A (n_3540), .B (n_3210), .C (n_3043), .D (n_1624), .Y(n_5538));
NOR2X1 g37500(.A (n_5290), .B (n_6594), .Y (n_4664));
NOR2X1 g37501(.A (n_5282), .B (n_6594), .Y (n_4663));
NAND2X1 g37502(.A (n_6972), .B (oc3_cfg_999), .Y (n_4662));
NAND4X1 g37051(.A (n_3106), .B (n_2943), .C (n_2473), .D (n_1506), .Y(n_5541));
AOI21X1 g37720(.A0 (n_5518), .A1 (n_1316), .B0 (n_2332), .Y (n_3919));
OAI21X1 g33618(.A0 (n_5030), .A1 (n_9286), .B0 (n_7924), .Y (n_9298));
OAI21X1 g33619(.A0 (n_5029), .A1 (n_9288), .B0 (n_7923), .Y (n_9297));
AOI21X1 g37721(.A0 (n_366), .A1 (n_2553), .B0 (n_2327), .Y (n_3918));
OAI21X1 g33614(.A0 (n_5034), .A1 (n_9307), .B0 (n_7930), .Y (n_9302));
OAI21X1 g33615(.A0 (n_5033), .A1 (n_9286), .B0 (n_7929), .Y (n_9301));
OAI21X1 g33616(.A0 (n_5032), .A1 (n_9235), .B0 (n_7927), .Y (n_9300));
OAI21X1 g33617(.A0 (n_5031), .A1 (n_9264), .B0 (n_7925), .Y (n_9299));
OAI21X1 g33610(.A0 (n_5040), .A1 (n_9286), .B0 (n_7935), .Y (n_9310));
OAI21X1 g33611(.A0 (n_5039), .A1 (n_9307), .B0 (n_7934), .Y (n_9308));
OAI21X1 g33613(.A0 (n_5035), .A1 (n_9307), .B0 (n_7932), .Y (n_9304));
NAND2X1 g34421(.A (u4_mem_b2_b_58 ), .B (n_7984), .Y (n_7995));
NAND2X1 g38911(.A (u3_mem_b3_b_139 ), .B (n_2463), .Y (n_2405));
NAND2X1 g37724(.A (n_2446), .B (n_2981), .Y (n_4600));
NAND2X1 g38914(.A (u4_mem_b3_b_130 ), .B (n_3546), .Y (n_3533));
NOR2X1 g41750(.A (n_465), .B (n_503), .Y (n_752));
AOI22X1 g37727(.A0 (n_6666), .A1 (n_2553), .B0 (n_6595), .B1(n_1316), .Y (n_2554));
XOR2X1 g35495(.A (n_5622), .B (n_4093), .Y (n_5623));
NAND2X1 g38889(.A (u6_mem_b3_b_146 ), .B (n_2465), .Y (n_2425));
AOI21X1 g38558(.A0 (u8_mem_b2_b_29 ), .A1 (n_4491), .B0 (n_2018), .Y(n_4278));
AOI21X1 g38559(.A0 (u8_mem_b1_b_63 ), .A1 (n_4502), .B0 (n_1930), .Y(n_4277));
AOI21X1 g38552(.A0 (u8_mem_b1_b_83 ), .A1 (n_4387), .B0 (n_2098), .Y(n_4281));
AOI21X1 g38553(.A0 (u8_mem_b1_b_85 ), .A1 (n_4387), .B0 (n_2009), .Y(n_4280));
AOI21X1 g38550(.A0 (u8_mem_b3_b_132 ), .A1 (n_3879), .B0 (n_1435), .Y(n_3841));
AOI21X1 g38551(.A0 (u8_mem_b1_b_81 ), .A1 (n_4387), .B0 (n_2036), .Y(n_4282));
AOI21X1 g38556(.A0 (u8_mem_b1_b_61 ), .A1 (n_4387), .B0 (n_2022), .Y(n_4279));
AOI21X1 g38557(.A0 (u3_mem_b1_b_70 ), .A1 (n_5148), .B0 (n_2698), .Y(n_4868));
AOI21X1 g38554(.A0 (u3_mem_b1_b ), .A1 (n_5148), .B0 (n_3412), .Y(n_4870));
AOI21X1 g38555(.A0 (u3_mem_b1_b_69 ), .A1 (n_5148), .B0 (n_2648), .Y(n_4869));
NAND2X1 g32626(.A (n_396), .B (n_9947), .Y (n_12019));
NAND2X1 g32624(.A (n_160), .B (n_10583), .Y (n_11632));
NAND2X1 g32625(.A (n_248), .B (n_9947), .Y (n_11985));
NAND2X1 g32622(.A (n_321), .B (n_9947), .Y (n_11989));
NAND2X1 g32623(.A (n_330), .B (n_9947), .Y (n_11675));
NAND2X1 g32620(.A (u11_wp_b3_b ), .B (n_9631), .Y (n_9834));
NAND2X1 g32621(.A (n_320), .B (n_9943), .Y (n_12009));
NAND2X1 g32628(.A (n_9514), .B (u9_wp_b3_b ), .Y (n_9686));
NAND2X1 g32629(.A (n_295), .B (n_9943), .Y (n_11949));
INVX1 g42750(.A (u6_wp_b2_b ), .Y (n_1255));
NAND2X1 g39091(.A (n_2465), .B (n_496), .Y (n_2360));
NAND2X1 g36679(.A (n_5255), .B (n_3966), .Y (n_5761));
OAI21X1 g36678(.A0 (n_4573), .A1 (n_5199), .B0 (n_784), .Y (n_6108));
OAI21X1 g36675(.A0 (n_12052), .A1 (n_12053), .B0 (n_784), .Y(n_6111));
OAI21X1 g36674(.A0 (n_12050), .A1 (n_12051), .B0 (n_784), .Y(n_6112));
OAI21X1 g36677(.A0 (n_5188), .A1 (n_5162), .B0 (n_634), .Y (n_5762));
OAI21X1 g36676(.A0 (n_12058), .A1 (n_12059), .B0 (n_784), .Y(n_6109));
OAI21X1 g36671(.A0 (n_12056), .A1 (n_12057), .B0 (n_784), .Y(n_6114));
OAI21X1 g36673(.A0 (n_12048), .A1 (n_12049), .B0 (n_784), .Y(n_6113));
NAND2X1 g45765(.A (n_12480), .B (n_12481), .Y (n_12482));
NAND4X1 g45767(.A (n_4114), .B (n_3098), .C (n_2291), .D (n_1383), .Y(n_12481));
NOR2X1 g45766(.A (u7_rp_b0_b ), .B (n_12640), .Y (n_12480));
OAI21X1 g45761(.A0 (n_5459), .A1 (n_5211), .B0 (n_12478), .Y(n_12479));
INVX1 g41376(.A (n_12682), .Y (n_3255));
INVX8 g41473(.A (n_1388), .Y (n_3117));
NOR2X1 g45762(.A (n_12640), .B (n_12634), .Y (n_12478));
NOR2X1 g30709(.A (n_10776), .B (n_12589), .Y (n_10963));
NOR2X1 g30708(.A (n_10825), .B (n_11128), .Y (n_11009));
AOI21X1 g30707(.A0 (n_415), .A1 (n_416), .B0 (n_9521), .Y (n_9617));
MX2X1 g40429(.A (crac_din_694), .B (in_slt_833), .S0 (n_1036), .Y(n_1047));
INVX1 g42341(.A (u11_mem_b2_b_116 ), .Y (n_125));
INVX1 g41422(.A (n_12803), .Y (n_1208));
INVX1 g41421(.A (n_1208), .Y (n_1391));
INVX2 g41427(.A (n_12747), .Y (n_4258));
NOR2X1 g41425(.A (n_564), .B (n_802), .Y (n_565));
MX2X1 g36019(.A (n_6514), .B (n_6604), .S0 (n_6649), .Y (n_6605));
MX2X1 g36018(.A (n_6607), .B (n_6563), .S0 (n_5341), .Y (n_6608));
MX2X1 g36011(.A (n_6646), .B (n_6620), .S0 (n_6908), .Y (n_6621));
MX2X1 g36010(.A (n_6623), .B (n_6570), .S0 (n_5341), .Y (n_6624));
MX2X1 g36013(.A (n_6539), .B (n_6614), .S0 (n_6908), .Y (n_6615));
MX2X1 g36012(.A (n_6618), .B (n_6617), .S0 (n_6908), .Y (n_6619));
MX2X1 g36014(.A (n_6883), .B (n_6922), .S0 (n_6908), .Y (n_6923));
MX2X1 g36017(.A (n_6610), .B (n_6602), .S0 (n_931), .Y (n_6611));
MX2X1 g36016(.A (n_6920), .B (n_6919), .S0 (n_6908), .Y (n_6921));
INVX1 g42311(.A (u9_mem_b3_b_58 ), .Y (n_6915));
INVX1 g42019(.A (u11_mem_b1_b_127 ), .Y (n_5984));
NAND2X1 g36901(.A (n_2547), .B (n_1239), .Y (n_4816));
NAND4X1 g36900(.A (n_4118), .B (n_2321), .C (n_3029), .D (n_1362), .Y(n_6264));
NOR2X1 g41373(.A (u13_ints_r_b25_b ), .B (n_608), .Y (n_609));
INVX1 g42472(.A (oc2_cfg_989), .Y (n_524));
INVX1 g34884(.A (n_9711), .Y (n_9688));
OR2X1 g34885(.A (u15_valid_r), .B (n_11827), .Y (n_9711));
NAND3X1 g34886(.A (n_7496), .B (n_2175), .C (n_9833), .Y (n_8676));
NAND2X1 g34731(.A (u7_mem_b1_b_82 ), .B (n_7651), .Y (n_7703));
NAND2X1 g34736(.A (u7_mem_b1_b_86 ), .B (n_7651), .Y (n_7698));
NAND2X1 g34737(.A (u8_mem_b2_b_54 ), .B (n_7976), .Y (n_7697));
NAND2X1 g34734(.A (u8_mem_b2_b_50 ), .B (n_7976), .Y (n_7700));
NAND2X1 g34735(.A (u7_mem_b1_b_85 ), .B (n_7651), .Y (n_7699));
NAND2X1 g34738(.A (u7_mem_b1_b_87 ), .B (n_7651), .Y (n_7696));
NOR2X1 g34888(.A (o4_status), .B (o4_status_972), .Y (n_7289));
NOR2X1 g34889(.A (o6_status), .B (o6_status_982), .Y (n_7288));
NOR2X1 g35281(.A (n_838), .B (rf_we), .Y (n_7287));
NAND3X1 g35280(.A (n_6330), .B (n_7011), .C (n_1460), .Y (n_7367));
NOR2X1 g35283(.A (n_7142), .B (n_11597), .Y (n_7366));
NOR2X1 g35282(.A (rf_we), .B (n_1300), .Y (n_7444));
INVX1 g35285(.A (n_8210), .Y (n_9359));
NOR2X1 g35284(.A (rf_we), .B (wb_addr_i_b4_b), .Y (n_7442));
NOR2X1 g35287(.A (n_7477), .B (n_1119), .Y (n_7481));
INVX1 g35286(.A (n_7481), .Y (n_8210));
NAND3X1 g35289(.A (n_5944), .B (n_6757), .C (n_2298), .Y (n_7285));
NOR2X1 g35288(.A (n_2574), .B (rf_we), .Y (n_7286));
OAI21X1 g35939(.A0 (n_5531), .A1 (n_7063), .B0 (n_6169), .Y (n_7060));
NAND2X1 g39277(.A (u4_mem_b2_b_53 ), .B (n_12087), .Y (n_3328));
NAND2X1 g39902(.A (u8_mem_b1_b_70 ), .B (n_12295), .Y (n_11460));
NAND2X1 g39903(.A (u8_mem_b2_b_52 ), .B (n_3441), .Y (n_2891));
NAND2X1 g39272(.A (u3_mem_b2_b_55 ), .B (n_3330), .Y (n_3331));
NAND2X1 g39901(.A (u8_mem_b1_b_85 ), .B (n_12291), .Y (n_3862));
MX2X1 g34088(.A (u7_mem_b0_b_103 ), .B (n_3647), .S0 (n_7493), .Y(n_9401));
MX2X1 g34089(.A (u7_mem_b0_b_104 ), .B (n_3684), .S0 (n_7493), .Y(n_9400));
MX2X1 g34084(.A (u7_mem_b0_b ), .B (n_3710), .S0 (n_7493), .Y(n_8753));
MX2X1 g34085(.A (u7_mem_b0_b_100 ), .B (n_3677), .S0 (n_7493), .Y(n_8752));
MX2X1 g34086(.A (u7_mem_b0_b_101 ), .B (n_3806), .S0 (n_7493), .Y(n_8751));
MX2X1 g34087(.A (u7_mem_b0_b_102 ), .B (n_3786), .S0 (n_7493), .Y(n_8750));
NAND2X1 g36939(.A (n_1646), .B (n_1640), .Y (n_4022));
AOI22X1 g40420(.A0 (u13_intm_r_b13_b ), .A1 (u13_ints_r_b13_b ), .B0(u13_intm_r_b15_b ), .B1 (u13_ints_r_b15_b ), .Y (n_557));
INVX1 g42010(.A (u11_mem_b3_b_85 ), .Y (n_5524));
INVX1 g42319(.A (u11_mem_b0_b_168 ), .Y (n_312));
AOI21X1 g35425(.A0 (n_6958), .A1 (n_4689), .B0 (n_7353), .Y (n_7348));
AOI21X1 g35424(.A0 (n_6971), .A1 (n_4735), .B0 (n_7353), .Y (n_7349));
AOI21X1 g35427(.A0 (n_6967), .A1 (n_4712), .B0 (n_7353), .Y (n_7346));
AOI21X1 g35426(.A0 (n_6968), .A1 (n_4715), .B0 (n_7353), .Y (n_7347));
AOI21X1 g35421(.A0 (n_6974), .A1 (n_4742), .B0 (n_7353), .Y (n_7352));
AOI21X1 g35420(.A0 (n_6969), .A1 (n_4693), .B0 (n_7353), .Y (n_7354));
AOI21X1 g35423(.A0 (n_6960), .A1 (n_4737), .B0 (n_7353), .Y (n_7350));
AOI21X1 g35422(.A0 (n_6973), .A1 (n_4692), .B0 (n_7353), .Y (n_7351));
AOI21X1 g35429(.A0 (n_6965), .A1 (n_4704), .B0 (n_7353), .Y (n_7344));
AOI21X1 g35428(.A0 (n_6966), .A1 (n_4709), .B0 (n_7353), .Y (n_7345));
INVX1 g42116(.A (u9_mem_b1_b_129 ), .Y (n_6551));
MX2X1 g40422(.A (crac_din_698), .B (in_slt_837), .S0 (n_1036), .Y(n_1022));
INVX4 g32817(.A (n_9741), .Y (n_10250));
INVX4 g32816(.A (n_10073), .Y (n_9741));
INVX4 g32811(.A (n_9741), .Y (n_10235));
MX2X1 g40425(.A (crac_din_702), .B (in_slt_841), .S0 (n_1036), .Y(n_1029));
INVX1 g43111(.A (u10_mem_b3_b_70 ), .Y (n_6588));
INVX1 g45357(.A (ic0_cfg), .Y (n_11578));
MX2X1 g40424(.A (crac_din_700), .B (in_slt_839), .S0 (n_1036), .Y(n_1028));
NOR2X1 g40072(.A (n_2864), .B (n_1985), .Y (n_2159));
NOR2X1 g40073(.A (n_2784), .B (n_2755), .Y (n_2785));
NOR2X1 g40070(.A (n_2712), .B (n_1985), .Y (n_2160));
NOR2X1 g40071(.A (n_1147), .B (n_2786), .Y (n_2787));
NOR2X1 g40076(.A (n_2831), .B (n_2057), .Y (n_2156));
NOR2X1 g40077(.A (n_2780), .B (n_2772), .Y (n_2781));
NAND2X1 g40074(.A (n_5157), .B (n_4533), .Y (n_2157));
NOR2X1 g40075(.A (n_2721), .B (n_2782), .Y (n_2783));
NOR2X1 g40078(.A (n_1082), .B (n_2786), .Y (n_2779));
NOR2X1 g40079(.A (n_2154), .B (n_2684), .Y (n_2155));
MX2X1 g40427(.A (crac_din_693), .B (in_slt_832), .S0 (n_1036), .Y(n_1194));
OAI21X1 g33529(.A0 (n_4451), .A1 (n_8333), .B0 (n_8028), .Y (n_8315));
AOI21X1 g37264(.A0 (n_5494), .A1 (n_6649), .B0 (n_4638), .Y (n_5495));
MX2X1 g37267(.A (u10_mem_b2_b_114 ), .B (n_4759), .S0 (n_5341), .Y(n_4760));
AOI21X1 g37266(.A0 (n_5490), .A1 (n_6649), .B0 (n_4651), .Y (n_5491));
AOI21X1 g37261(.A0 (n_5498), .A1 (n_6649), .B0 (n_4650), .Y (n_5499));
MX2X1 g37260(.A (u10_mem_b2_b_113 ), .B (n_4761), .S0 (n_5341), .Y(n_4762));
MX2X1 g37263(.A (u10_mem_b1_b_149 ), .B (n_5339), .S0 (n_6475), .Y(n_5349));
AOI21X1 g37262(.A0 (n_5496), .A1 (n_6649), .B0 (n_4637), .Y (n_5497));
MX2X1 g37269(.A (u9_mem_b2_b_112 ), .B (n_4755), .S0 (n_5732), .Y(n_4756));
MX2X1 g37268(.A (u9_mem_b2_b_110 ), .B (n_4757), .S0 (n_6898), .Y(n_4758));
NOR2X1 g41211(.A (u13_ints_r_b13_b ), .B (n_490), .Y (n_597));
NAND2X1 g41210(.A (n_5225), .B (n_1300), .Y (n_7019));
INVX1 g41213(.A (n_6042), .Y (n_1200));
OR2X1 g41212(.A (n_1301), .B (n_5831), .Y (n_1302));
NOR2X1 g41215(.A (u13_ints_r_b4_b ), .B (n_492), .Y (n_733));
AND2X1 g41214(.A (n_838), .B (wb_addr_i_b3_b), .Y (n_6042));
NOR2X1 g41217(.A (n_598), .B (n_804), .Y (n_599));
OR2X1 g41216(.A (n_7017), .B (n_12585), .Y (n_1146));
NOR2X1 g41219(.A (n_699), .B (n_872), .Y (n_700));
OAI21X1 g31049(.A0 (n_5299), .A1 (n_10820), .B0 (n_10361), .Y(n_10862));
OAI21X1 g31048(.A0 (n_5305), .A1 (n_10880), .B0 (n_10362), .Y(n_10863));
AOI22X1 g31739(.A0 (n_7447), .A1 (n_7528), .B0 (n_569), .B1 (n_7378),.Y (n_8909));
AOI22X1 g31738(.A0 (n_7449), .A1 (n_7531), .B0 (n_700), .B1 (n_7379),.Y (n_8915));
NAND3X1 g31735(.A (n_12531), .B (n_12149), .C (n_991), .Y (n_10954));
AOI21X1 g31734(.A0 (n_2986), .A1 (n_4836), .B0 (n_12339), .Y(n_9973));
OAI21X1 g31041(.A0 (n_5314), .A1 (n_10820), .B0 (n_10367), .Y(n_10870));
NAND3X1 g31736(.A (n_1229), .B (n_12608), .C (n_9833), .Y (n_10950));
OAI21X1 g31047(.A0 (n_5423), .A1 (n_10450), .B0 (n_9987), .Y(n_10675));
OAI21X1 g31046(.A0 (n_5308), .A1 (n_10820), .B0 (n_10363), .Y(n_10864));
AND2X1 g31732(.A (n_5625), .B (ac97_rst_force), .Y (n_9492));
AOI22X1 g33399(.A0 (n_4389), .A1 (n_7505), .B0 (n_7758), .B1(u6_wp_b2_b ), .Y (n_8477));
AOI22X1 g33398(.A0 (n_4349), .A1 (n_7496), .B0 (n_7870), .B1(u5_wp_b2_b ), .Y (n_8478));
AOI22X1 g33395(.A0 (n_2487), .A1 (n_7490), .B0 (n_7976), .B1(u8_wp_b2_b ), .Y (n_8481));
OR2X1 g33394(.A (n_5439), .B (n_7519), .Y (n_7520));
AOI22X1 g33397(.A0 (n_4395), .A1 (n_7499), .B0 (n_7984), .B1(u4_wp_b2_b ), .Y (n_8479));
AOI22X1 g33396(.A0 (n_4333), .A1 (n_7423), .B0 (n_8101), .B1(u3_wp_b2_b ), .Y (n_8480));
AOI21X1 g33391(.A0 (n_1120), .A1 (n_7478), .B0 (n_1289), .Y (n_8482));
AOI21X1 g33390(.A0 (n_1126), .A1 (n_7479), .B0 (n_1259), .Y (n_8483));
OR2X1 g33393(.A (n_5596), .B (n_7446), .Y (n_7447));
OR2X1 g33392(.A (n_5597), .B (n_7448), .Y (n_7449));
MX2X1 g34000(.A (u4_mem_b0_b_117 ), .B (n_3764), .S0 (n_7499), .Y(n_8821));
INVX1 g42776(.A (u9_mem_b3_b_63 ), .Y (n_6909));
NAND2X1 g39234(.A (u5_mem_b2_b_33 ), .B (n_12823), .Y (n_12810));
INVX1 g42770(.A (u9_mem_b2_b_108 ), .Y (n_35));
INVX1 g42746(.A (n_12581), .Y (n_771));
NAND2X1 g37579(.A (n_5480), .B (n_3060), .Y (n_4639));
INVX1 g42745(.A (n_771), .Y (n_886));
INVX1 g42742(.A (u10_mem_b0_b_160 ), .Y (n_6384));
INVX2 g42741(.A (oc1_cfg), .Y (n_458));
INVX1 g42173(.A (u9_mem_b2_b_101 ), .Y (n_6638));
NOR2X1 g39236(.A (n_3117), .B (n_2763), .Y (n_3346));
NAND2X1 g39599(.A (u4_mem_b2_b_29 ), .B (n_12087), .Y (n_2277));
AOI21X1 g35639(.A0 (n_6325), .A1 (n_5756), .B0 (n_7214), .Y (n_7227));
AOI21X1 g35630(.A0 (n_6296), .A1 (n_6099), .B0 (n_12640), .Y(n_7235));
AOI21X1 g35631(.A0 (n_6295), .A1 (n_6097), .B0 (n_12640), .Y(n_7233));
AOI21X1 g35632(.A0 (n_6308), .A1 (n_6096), .B0 (n_12640), .Y(n_7232));
NAND2X1 g39595(.A (n_12369), .B (u6_mem_b0_b_116 ), .Y (n_3073));
NAND2X1 g39594(.A (u6_mem_b1_b_85 ), .B (n_4253), .Y (n_4163));
AOI21X1 g35636(.A0 (n_6293), .A1 (n_6095), .B0 (n_12640), .Y(n_7230));
AOI21X1 g35637(.A0 (n_5914), .A1 (n_6761), .B0 (n_12640), .Y(n_7306));
NAND4X1 g37576(.A (n_1051), .B (n_449), .C (n_742), .D (u2_to_cnt_b0_b), .Y (n_5629));
AOI22X1 g38783(.A0 (n_3316), .A1 (n_634), .B0 (n_6316), .B1 (n_763),.Y (n_4267));
INVX1 g42453(.A (n_403), .Y (n_1206));
NAND2X1 g41172(.A (u4_rp_b2_b ), .B (n_551), .Y (n_552));
OAI21X1 g38782(.A0 (n_12262), .A1 (n_145), .B0 (n_929), .Y (n_4268));
INVX1 g42568(.A (u11_mem_b0_b_174 ), .Y (n_1610));
INVX2 g41173(.A (n_5876), .Y (n_7115));
NAND2X1 g37573(.A (n_5645), .B (n_4206), .Y (n_5228));
AND2X1 g41174(.A (oc2_cfg_985), .B (n_242), .Y (n_5876));
OR2X1 g37572(.A (n_1777), .B (ac97_reset_pad_o_), .Y (n_1778));
INVX1 g42296(.A (u11_mem_b2_b_102 ), .Y (n_6460));
INVX1 g31767(.A (n_9606), .Y (n_9607));
NAND2X1 g39735(.A (n_12839), .B (u4_mem_b0_b_96 ), .Y (n_12829));
NAND2X1 g39042(.A (u8_mem_b2_b_55 ), .B (n_2366), .Y (n_2367));
NAND2X1 g39041(.A (u3_mem_b2_b_53 ), .B (n_3330), .Y (n_2640));
NAND2X1 g39040(.A (in_slt_406), .B (n_4623), .Y (n_4239));
NAND2X1 g39047(.A (n_4560), .B (in_slt_451), .Y (n_5313));
INVX1 g39046(.A (n_5313), .Y (n_4237));
NAND2X1 g39045(.A (n_4560), .B (in_slt_448), .Y (n_5335));
INVX1 g39044(.A (n_5335), .Y (n_4238));
NAND2X1 g39049(.A (u3_mem_b1_b_77 ), .B (n_3316), .Y (n_3489));
NAND2X1 g39048(.A (n_12839), .B (u4_mem_b0_b_117 ), .Y (n_3490));
NAND2X1 g39739(.A (u4_mem_b1_b_66 ), .B (n_12273), .Y (n_11659));
NOR2X1 g39738(.A (n_3332), .B (n_2829), .Y (n_2987));
NAND2X1 g36811(.A (n_1694), .B (n_1693), .Y (n_4041));
NAND2X1 g36810(.A (n_1674), .B (n_1710), .Y (n_4042));
NAND2X1 g36813(.A (n_1709), .B (n_1696), .Y (n_4040));
OR2X1 g36812(.A (n_1815), .B (wb_we_i), .Y (n_1814));
NAND2X1 g36815(.A (n_1702), .B (n_1731), .Y (n_4039));
NAND2X1 g36814(.A (n_1862), .B (n_3893), .Y (n_4824));
NAND4X1 g36817(.A (n_12829), .B (n_12830), .C (n_2849), .D (n_3534),.Y (n_6252));
INVX1 g36816(.A (n_6252), .Y (n_5729));
NAND4X1 g36819(.A (n_11445), .B (n_11446), .C (n_2363), .D (n_2393),.Y (n_5798));
INVX1 g36818(.A (n_5798), .Y (n_5572));
INVX1 g43010(.A (u10_mem_b0_b_153 ), .Y (n_6337));
NAND2X1 g39115(.A (n_3339), .B (in_slt_429), .Y (n_5282));
NOR2X1 g40275(.A (n_2103), .B (n_2829), .Y (n_1994));
NOR2X1 g40276(.A (n_2755), .B (n_1985), .Y (n_1993));
NAND2X1 g39116(.A (n_12369), .B (u6_mem_b0_b_115 ), .Y (n_3437));
NOR2X1 g40270(.A (n_2038), .B (n_2765), .Y (n_1997));
NOR2X1 g40271(.A (n_2689), .B (n_2712), .Y (n_2690));
NAND2X1 g39890(.A (n_12839), .B (u4_mem_b0_b_106 ), .Y (n_12827));
NOR2X1 g40272(.A (n_2705), .B (n_2686), .Y (n_2688));
NOR2X1 g40273(.A (n_2093), .B (n_2707), .Y (n_1996));
NAND2X1 g39892(.A (u3_mem_b2_b_46 ), .B (n_12619), .Y (n_2898));
OR2X1 g41423_dup(.A (n_524), .B (n_447), .Y (n_12804));
OAI21X1 g35861(.A0 (n_5727), .A1 (n_11934), .B0 (n_6778), .Y(n_7199));
INVX1 g39895(.A (n_4747), .Y (n_2895));
INVX1 g41989(.A (u9_mem_b1_b_128 ), .Y (n_6656));
AOI21X1 g38303(.A0 (u5_mem_b2_b ), .A1 (n_4378), .B0 (n_2210), .Y(n_4379));
AOI21X1 g35647(.A0 (n_5910), .A1 (n_5745), .B0 (n_7120), .Y (n_7123));
AOI21X1 g38302(.A0 (u8_mem_b1_b_75 ), .A1 (n_4387), .B0 (n_2215), .Y(n_4380));
INVX1 g41981(.A (u10_mem_b3_b_59 ), .Y (n_6575));
AND2X1 g40278(.A (n_476), .B (n_869), .Y (n_870));
INVX1 g41983(.A (n_4734), .Y (n_568));
NAND2X1 g39549(.A (u7_mem_b2_b_39 ), .B (n_12654), .Y (n_3098));
NAND2X1 g37173(.A (n_2511), .B (n_2359), .Y (n_6008));
NOR2X1 g40279(.A (n_935), .B (n_2792), .Y (n_1991));
NAND2X1 g39898(.A (n_12825), .B (u3_mem_b0_b_109 ), .Y (n_2894));
AOI21X1 g38300(.A0 (u6_mem_b1_b_85 ), .A1 (n_5112), .B0 (n_2668), .Y(n_5011));
NAND2X1 g39547(.A (u8_mem_b1_b_74 ), .B (n_12295), .Y (n_11462));
AOI21X1 g38307(.A0 (u5_mem_b2_b_40 ), .A1 (n_4378), .B0 (n_2221), .Y(n_4375));
NAND2X1 g39544(.A (n_2491), .B (u7_mem_b0_b_113 ), .Y (n_1807));
AOI21X1 g38306(.A0 (u5_mem_b2_b_39 ), .A1 (n_4378), .B0 (n_2007), .Y(n_4376));
NAND2X1 g39545(.A (n_12204), .B (u6_mem_b0_b ), .Y (n_11751));
NAND2X1 g37177(.A (n_3895), .B (n_2329), .Y (n_6444));
NOR2X1 g39542(.A (n_3453), .B (n_2790), .Y (n_3103));
NAND2X1 g37176(.A (n_2517), .B (n_2922), .Y (n_5993));
INVX1 g42234(.A (u11_mem_b2_b_104 ), .Y (n_5978));
NAND2X1 g39543(.A (u8_mem_b1_b_60 ), .B (n_12295), .Y (n_11499));
OAI21X1 g33553(.A0 (n_4427), .A1 (n_9346), .B0 (n_8004), .Y (n_8285));
OAI21X1 g33552(.A0 (n_4428), .A1 (n_9333), .B0 (n_8005), .Y (n_8286));
OAI21X1 g33551(.A0 (n_4327), .A1 (n_8318), .B0 (n_8006), .Y (n_8287));
OAI21X1 g33550(.A0 (n_4429), .A1 (n_8333), .B0 (n_8007), .Y (n_8289));
OAI21X1 g33557(.A0 (n_4422), .A1 (n_9326), .B0 (n_8000), .Y (n_8281));
NAND2X1 g34276(.A (u8_mem_b1_b_62 ), .B (n_7976), .Y (n_8124));
OAI21X1 g33803(.A0 (n_5115), .A1 (n_9022), .B0 (n_8077), .Y (n_9069));
OAI21X1 g33554(.A0 (n_4426), .A1 (n_8333), .B0 (n_8003), .Y (n_8284));
OAI21X1 g33559(.A0 (n_4420), .A1 (n_8333), .B0 (n_7998), .Y (n_8278));
OAI21X1 g33558(.A0 (n_4421), .A1 (n_8333), .B0 (n_7999), .Y (n_8280));
OAI21X1 g33809(.A0 (n_4858), .A1 (n_8856), .B0 (n_7568), .Y (n_9063));
OAI21X1 g33808(.A0 (n_4918), .A1 (n_9055), .B0 (n_7719), .Y (n_9064));
INVX1 g42235(.A (u10_mem_b1_b ), .Y (n_5981));
INVX1 g37078(.A (n_6172), .Y (n_5679));
NAND4X1 g37079(.A (n_11729), .B (n_11730), .C (n_2872), .D (n_1518),.Y (n_6172));
INVX1 g37070(.A (n_12618), .Y (n_5682));
MX2X1 g38711(.A (u7_mem_b0_b_121 ), .B (wb_din_691), .S0 (n_3622), .Y(n_3635));
NOR2X1 g37072(.A (n_3875), .B (n_2368), .Y (n_4805));
NAND2X1 g37073(.A (n_2503), .B (n_1707), .Y (n_3999));
MX2X1 g38714(.A (u6_mem_b0_b_91 ), .B (wb_din_661), .S0 (n_3632), .Y(n_3630));
MX2X1 g38715(.A (u6_mem_b0_b_93 ), .B (wb_din_663), .S0 (n_3632), .Y(n_3628));
MX2X1 g38717(.A (u7_mem_b0_b_99 ), .B (wb_din_669), .S0 (n_3622), .Y(n_3626));
AOI21X1 g38504(.A0 (u7_mem_b2_b_59 ), .A1 (n_4509), .B0 (n_2026), .Y(n_4307));
INVX1 g42233(.A (u10_mem_b0_b_161 ), .Y (n_6382));
NAND2X1 g38809(.A (u8_mem_b3_b_147 ), .B (n_2468), .Y (n_1812));
INVX2 g42765(.A (ic0_cfg_1025), .Y (n_836));
NAND2X1 g38879(.A (u3_mem_b3_b_143 ), .B (n_2463), .Y (n_2432));
NAND2X1 g32607(.A (n_9453), .B (oc0_int_set_708), .Y (n_9578));
NAND2X1 g32608(.A (n_9452), .B (oc1_int_set_710), .Y (n_9577));
NAND2X1 g32609(.A (n_9451), .B (oc2_int_set_712), .Y (n_9576));
NOR2X1 g35572(.A (n_1085), .B (i3_re), .Y (n_6713));
OAI21X1 g36657(.A0 (n_3915), .A1 (n_4596), .B0 (n_5772), .Y (n_5773));
OAI21X1 g36656(.A0 (n_4570), .A1 (n_4597), .B0 (n_5772), .Y (n_5774));
OAI21X1 g36655(.A0 (n_3916), .A1 (n_4598), .B0 (n_6091), .Y (n_5775));
OAI21X1 g36654(.A0 (n_3917), .A1 (n_4599), .B0 (n_6091), .Y (n_5776));
NAND2X1 g36653(.A (n_5251), .B (n_2614), .Y (n_5777));
NAND2X1 g36651(.A (n_5256), .B (n_3969), .Y (n_5779));
OAI21X1 g36659(.A0 (n_4593), .A1 (n_4592), .B0 (n_5772), .Y (n_5770));
OAI21X1 g36658(.A0 (n_3914), .A1 (n_4594), .B0 (n_5772), .Y (n_5771));
NAND2X1 g36389(.A (n_6150), .B (n_6316), .Y (n_11987));
NAND2X1 g36388(.A (n_5813), .B (n_2567), .Y (n_5910));
AND2X1 g45744(.A (n_634), .B (n_12535), .Y (n_12457));
OAI21X1 g45743(.A0 (n_5186), .A1 (n_5187), .B0 (n_12457), .Y(n_12458));
NAND2X1 g45742(.A (n_12458), .B (n_12459), .Y (n_12460));
OAI21X1 g45741(.A0 (n_5680), .A1 (n_7077), .B0 (n_6188), .Y(n_12454));
NAND2X1 g38870(.A (u4_mem_b3_b_145 ), .B (n_3556), .Y (n_3537));
NAND2X1 g36381(.A (n_12618), .B (n_6316), .Y (n_6289));
NAND2X1 g36380(.A (n_6235), .B (n_6316), .Y (n_6290));
NAND2X1 g36382(.A (n_12755), .B (n_6316), .Y (n_6288));
NAND2X1 g36385(.A (n_5798), .B (n_2567), .Y (n_5911));
NAND2X1 g36384(.A (n_12116), .B (n_6316), .Y (n_6287));
NAND2X1 g36387(.A (n_6260), .B (n_2567), .Y (n_6286));
NAND2X1 g36386(.A (n_11925), .B (n_6824), .Y (n_6818));
NAND2X1 g38872(.A (u7_mem_b3_b_143 ), .B (n_1546), .Y (n_1339));
NAND2X1 g38875(.A (u7_mem_b3_b_152 ), .B (n_1546), .Y (n_1536));
NAND2X1 g38874(.A (u7_mem_b3_b_134 ), .B (n_1538), .Y (n_1537));
OAI21X1 g37382(.A0 (u9_mem_b0_b_172 ), .A1 (n_6856), .B0 (n_4672), .Y(n_5483));
OAI21X1 g37380(.A0 (u9_mem_b0_b_169 ), .A1 (n_6856), .B0 (n_4646), .Y(n_5486));
OAI21X1 g37386(.A0 (u9_mem_b0_b_176 ), .A1 (n_6856), .B0 (n_4667), .Y(n_5477));
OAI21X1 g37387(.A0 (u9_mem_b0_b_177 ), .A1 (n_6856), .B0 (n_4669), .Y(n_5475));
OAI21X1 g37385(.A0 (u9_mem_b0_b_175 ), .A1 (n_6856), .B0 (n_4671), .Y(n_5479));
OAI21X1 g37388(.A0 (u9_mem_b0_b_178 ), .A1 (n_6856), .B0 (n_4668), .Y(n_5474));
OAI21X1 g37389(.A0 (u9_mem_b0_b_179 ), .A1 (n_6856), .B0 (n_4670), .Y(n_5473));
AOI21X1 g38578(.A0 (u3_mem_b1_b_85 ), .A1 (n_5148), .B0 (n_2704), .Y(n_4856));
AOI21X1 g38579(.A0 (u3_mem_b1_b_86 ), .A1 (n_5157), .B0 (n_2723), .Y(n_4855));
MX2X1 g36033(.A (n_6014), .B (n_6013), .S0 (n_6594), .Y (n_6015));
MX2X1 g36032(.A (n_6586), .B (n_6585), .S0 (n_6594), .Y (n_6587));
MX2X1 g36031(.A (n_6589), .B (n_6588), .S0 (n_6594), .Y (n_6590));
MX2X1 g36030(.A (n_6592), .B (n_6591), .S0 (n_6594), .Y (n_6593));
MX2X1 g36037(.A (n_5997), .B (n_6005), .S0 (n_6594), .Y (n_6006));
MX2X1 g36036(.A (n_6008), .B (n_6007), .S0 (n_6594), .Y (n_6009));
MX2X1 g36035(.A (n_6900), .B (n_6899), .S0 (n_6898), .Y (n_6901));
MX2X1 g36034(.A (n_6011), .B (n_6010), .S0 (n_6594), .Y (n_6012));
MX2X1 g36039(.A (n_6579), .B (n_6578), .S0 (n_6594), .Y (n_6580));
MX2X1 g36038(.A (n_6582), .B (n_6581), .S0 (n_6908), .Y (n_6583));
INVX1 g42842(.A (u3_wp_b1_b ), .Y (n_626));
NAND2X1 g39530(.A (u7_mem_b2_b_50 ), .B (n_12645), .Y (n_4175));
NOR2X1 g40318(.A (n_2083), .B (n_2707), .Y (n_1963));
NOR2X1 g37042(.A (u26_ps_cnt_b3_b ), .B (n_818), .Y (n_1014));
NAND2X1 g39452(.A (u5_mem_b1_b_62 ), .B (n_3236), .Y (n_11440));
NOR2X1 g39537(.A (n_2767), .B (n_1488), .Y (n_1283));
NAND2X1 g39310(.A (u5_mem_b1_b_79 ), .B (n_3236), .Y (n_3288));
MX2X1 g31384(.A (u11_din_tmp_48), .B (in_slt_451), .S0 (n_10103), .Y(n_10098));
MX2X1 g31385(.A (u11_din_tmp_49), .B (in_slt_452), .S0 (n_10103), .Y(n_10097));
MX2X1 g31386(.A (u11_din_tmp_50), .B (in_slt_453), .S0 (n_10103), .Y(n_10096));
MX2X1 g31387(.A (u10_din_tmp1), .B (in_slt_422), .S0 (n_9860), .Y(n_9861));
MX2X1 g31380(.A (u11_din_tmp_44), .B (in_slt_447), .S0 (n_10103), .Y(n_10102));
MX2X1 g31381(.A (u11_din_tmp_45), .B (in_slt_448), .S0 (n_10103), .Y(n_10101));
MX2X1 g31382(.A (u11_din_tmp_46), .B (in_slt_449), .S0 (n_10103), .Y(n_10100));
MX2X1 g31383(.A (u11_din_tmp_47), .B (in_slt_450), .S0 (n_10103), .Y(n_10099));
MX2X1 g31388(.A (u10_din_tmp_51), .B (in_slt_432), .S0 (n_9860), .Y(n_9859));
MX2X1 g31389(.A (u10_din_tmp_52), .B (in_slt_433), .S0 (n_9860), .Y(n_9858));
NOR2X1 g39453(.A (n_3332), .B (n_2792), .Y (n_3169));
NAND2X1 g37927(.A (n_4124), .B (n_2479), .Y (n_5457));
NAND2X1 g37924(.A (n_1535), .B (n_4142), .Y (n_5459));
NAND2X1 g37925(.A (n_4223), .B (n_2952), .Y (n_5458));
NAND2X1 g37922(.A (n_4214), .B (n_3389), .Y (n_5460));
NAND2X1 g37920(.A (n_1547), .B (n_4126), .Y (n_5461));
AOI22X1 g37921(.A0 (n_4097), .A1 (in_slt_451), .B0 (n_2325), .B1(in_slt_449), .Y (n_3894));
NAND2X1 g37128(.A (n_1865), .B (n_1663), .Y (n_3998));
NAND2X1 g37928(.A (n_4203), .B (n_3253), .Y (n_5456));
AOI22X1 g37929(.A0 (u10_din_tmp_44), .A1 (n_3339), .B0 (n_3911), .B1(in_slt_423), .Y (n_4558));
AND2X1 g41404(.A (wb_we_i), .B (wb_stb_i), .Y (n_869));
NAND2X1 g39090(.A (n_1546), .B (n_457), .Y (n_1500));
NOR2X1 g41406(.A (n_175), .B (n_571), .Y (n_683));
INVX1 g41155(.A (n_1409), .Y (n_2696));
BUFX3 g41152(.A (n_1147), .Y (n_5019));
INVX1 g41153(.A (n_1409), .Y (n_2689));
NAND2X1 g41150(.A (n_431), .B (n_4706), .Y (n_1148));
INVX1 g33231(.A (o9_empty), .Y (n_9532));
NOR2X1 g40314(.A (n_2020), .B (n_2684), .Y (n_1967));
AOI21X1 g38506(.A0 (u7_mem_b2_b_34 ), .A1 (n_4509), .B0 (n_1997), .Y(n_4305));
NAND2X1 g39760(.A (u8_mem_b1_b_76 ), .B (n_12295), .Y (n_11669));
NOR2X1 g39454(.A (n_3332), .B (n_2729), .Y (n_3167));
INVX1 g41159(.A (n_1409), .Y (n_2749));
INVX1 g42175(.A (u9_mem_b3_b_87 ), .Y (n_5350));
INVX1 g42174(.A (u10_mem_b3_b_69 ), .Y (n_6591));
NAND2X1 g39093(.A (n_2344), .B (in_slt_419), .Y (n_2359));
NAND2X1 g34718(.A (u7_mem_b1_b_70 ), .B (n_7651), .Y (n_7719));
NAND2X1 g34719(.A (u7_mem_b1_b_71 ), .B (n_7651), .Y (n_7718));
NAND2X1 g34868(.A (u8_mem_b2_b_55 ), .B (n_7976), .Y (n_7566));
NAND2X1 g34869(.A (u3_mem_b1_b_84 ), .B (n_8101), .Y (n_7565));
NAND2X1 g34866(.A (u3_mem_b1_b_82 ), .B (n_8101), .Y (n_7568));
NAND2X1 g34867(.A (u8_mem_b2_b_53 ), .B (n_7976), .Y (n_7567));
NAND2X1 g34716(.A (u7_mem_b1_b ), .B (n_7651), .Y (n_7722));
NAND2X1 g34717(.A (u7_mem_b1_b_69 ), .B (n_7651), .Y (n_7721));
NAND2X1 g34862(.A (u3_mem_b1_b_80 ), .B (n_8101), .Y (n_7572));
OR2X1 g34711(.A (i6_status), .B (n_7439), .Y (n_7440));
NAND2X1 g34860(.A (u8_mem_b2_b_46 ), .B (n_7976), .Y (n_7574));
NAND2X1 g34861(.A (u8_mem_b2_b_29 ), .B (n_7976), .Y (n_7573));
NAND2X1 g39096(.A (n_12204), .B (u6_mem_b0_b_105 ), .Y (n_11703));
NOR2X1 g31568(.A (n_9803), .B (n_6752), .Y (n_10399));
NAND2X1 g31569(.A (n_3992), .B (n_12589), .Y (n_11513));
AOI22X1 g37881(.A0 (u11_din_tmp_51), .A1 (n_4560), .B0 (n_4097), .B1(in_slt_452), .Y (n_3907));
NAND2X1 g39765(.A (u7_mem_b2_b ), .B (n_12641), .Y (n_2971));
NAND2X1 g39455(.A (u4_mem_b2_b_38 ), .B (n_12079), .Y (n_3166));
NAND2X1 g39534(.A (u4_mem_b2_b_51 ), .B (n_12091), .Y (n_3109));
NAND2X1 g39928(.A (u3_mem_b2_b_48 ), .B (n_3330), .Y (n_2870));
NAND2X1 g39929(.A (n_12840), .B (u4_mem_b0_b_99 ), .Y (n_11662));
NAND2X1 g39920(.A (u8_mem_b1_b_75 ), .B (n_12301), .Y (n_12037));
NAND2X1 g39921(.A (u6_mem_b1_b_63 ), .B (n_4253), .Y (n_11710));
NAND2X1 g39922(.A (u8_mem_b2_b_58 ), .B (n_3441), .Y (n_3866));
NAND2X1 g39923(.A (u3_mem_b1_b_64 ), .B (n_3316), .Y (n_2874));
NAND2X1 g39925(.A (u5_mem_b2_b_55 ), .B (n_12823), .Y (n_2235));
NAND2X1 g39926(.A (u3_mem_b2_b_32 ), .B (n_3207), .Y (n_2872));
NAND2X1 g39927(.A (u3_mem_b1_b_89 ), .B (n_3316), .Y (n_2871));
NAND2X1 g39559(.A (n_12204), .B (u6_mem_b0_b_97 ), .Y (n_11715));
OAI21X1 g37383(.A0 (u9_mem_b0_b_173 ), .A1 (n_5480), .B0 (n_4677), .Y(n_5482));
INVX1 g41988(.A (oc1_int_set_710), .Y (n_488));
NAND2X1 g39274(.A (n_2344), .B (in_slt_424), .Y (n_2334));
XOR2X1 g37202(.A (u26_ps_cnt_b4_b ), .B (n_1449), .Y (n_3994));
NAND2X1 g39275(.A (n_2491), .B (u7_mem_b0_b_107 ), .Y (n_2333));
XOR2X1 g40448(.A (u11_wp_b0_b ), .B (u11_wp_b1_b ), .Y (n_825));
XOR2X1 g40447(.A (u9_rp_b1_b ), .B (u9_wp_b2_b ), .Y (n_1188));
INVX1 g35406(.A (i3_status_1022), .Y (n_6718));
XOR2X1 g40445(.A (n_12634), .B (n_1921), .Y (n_4797));
XOR2X1 g40444(.A (n_9641), .B (u10_wp_b1_b ), .Y (n_1189));
XOR2X1 g40443(.A (n_1033), .B (n_3559), .Y (n_2594));
XOR2X1 g40442(.A (u10_rp_b1_b ), .B (u10_wp_b2_b ), .Y (n_786));
XOR2X1 g40441(.A (n_6821), .B (n_11585), .Y (n_4799));
XOR2X1 g40440(.A (n_1923), .B (n_6824), .Y (n_4801));
NAND2X1 g39555(.A (u6_mem_b1_b_74 ), .B (n_4253), .Y (n_11704));
OAI21X1 g45678(.A0 (n_12376), .A1 (n_11673), .B0 (n_12377), .Y(n_12378));
AND2X1 g32837(.A (n_12689), .B (n_12534), .Y (n_11136));
INVX1 g32836(.A (n_11136), .Y (n_9907));
NAND2X1 g32835(.A (n_3942), .B (n_9447), .Y (n_9572));
INVX2 g32834(.A (n_9572), .Y (n_9633));
OAI21X1 g37200(.A0 (u11_rp_b1_b ), .A1 (n_853), .B0 (n_1121), .Y(n_4081));
NOR2X1 g32839(.A (n_9362), .B (n_5839), .Y (n_9519));
NAND2X1 g39129(.A (n_12825), .B (u3_mem_b0_b_121 ), .Y (n_3429));
INVX1 g41864(.A (u9_mem_b2_b_100 ), .Y (n_6641));
NAND2X1 g39554(.A (u8_mem_b2_b_47 ), .B (n_2366), .Y (n_2287));
NAND2X1 g34355(.A (u4_mem_b1_b_74 ), .B (n_7984), .Y (n_8048));
NAND2X1 g40(.A (u4_mem_b2_b_41 ), .B (n_12079), .Y (n_12741));
NAND2X1 g41(.A (n_11897), .B (n_11900), .Y (n_11901));
NAND2X1 g42(.A (n_11895), .B (n_12115), .Y (n_11897));
NAND2X1 g43(.A (n_11898), .B (n_12664), .Y (n_11900));
NAND4X1 g44(.A (n_2874), .B (n_11737), .C (n_11738), .D (n_1507), .Y(n_11895));
NAND4X1 g45(.A (n_3701), .B (n_3150), .C (n_3383), .D (n_1511), .Y(n_11898));
NAND2X1 g48(.A (n_12634), .B (n_6202), .Y (n_12121));
OAI21X1 g49(.A0 (n_5683), .A1 (n_7077), .B0 (n_6220), .Y (n_11908));
NAND2X1 g31700(.A (n_96), .B (n_10081), .Y (n_9987));
OR2X1 g32976_dup(.A (n_12636), .B (n_12501), .Y (n_11890));
AOI22X1 g37796(.A0 (n_1756), .A1 (n_312), .B0 (n_1644), .B1 (n_1643),.Y (n_1645));
NOR2X1 g40058(.A (n_1147), .B (n_2792), .Y (n_2797));
NOR2X1 g40059(.A (n_867), .B (n_2786), .Y (n_2167));
NAND2X1 g39556(.A (u6_mem_b2_b_36 ), .B (n_2285), .Y (n_2286));
MX2X1 g38655(.A (u5_mem_b0_b_91 ), .B (wb_din_661), .S0 (n_3720), .Y(n_3724));
NOR2X1 g40056(.A (n_2784), .B (n_2804), .Y (n_2800));
NOR2X1 g40057(.A (n_2784), .B (n_2818), .Y (n_2799));
NOR2X1 g40050(.A (n_2765), .B (n_2182), .Y (n_2174));
NOR2X1 g40051(.A (n_2788), .B (n_3008), .Y (n_2803));
NOR2X1 g40052(.A (n_941), .B (n_2716), .Y (n_2173));
NOR2X1 g40053(.A (n_2770), .B (n_2801), .Y (n_2802));
AOI21X1 g38389(.A0 (u8_mem_b3_b_129 ), .A1 (n_3879), .B0 (n_1477), .Y(n_3857));
AOI21X1 g38383(.A0 (u3_mem_b2_b_47 ), .A1 (n_4533), .B0 (n_1938), .Y(n_4347));
AOI21X1 g38382(.A0 (u3_mem_b2_b_38 ), .A1 (n_4533), .B0 (n_2010), .Y(n_4348));
AOI21X1 g38381(.A0 (u7_mem_b3_b_148 ), .A1 (n_5145), .B0 (n_2879), .Y(n_4959));
AOI21X1 g38380(.A0 (u3_mem_b3_b_146 ), .A1 (n_5133), .B0 (n_3467), .Y(n_4960));
AOI21X1 g38387(.A0 (u7_mem_b3_b_125 ), .A1 (n_5145), .B0 (n_2907), .Y(n_4957));
AOI21X1 g38386(.A0 (u3_mem_b3_b_142 ), .A1 (n_5133), .B0 (n_2961), .Y(n_4958));
AOI21X1 g38385(.A0 (u3_mem_b2_b_48 ), .A1 (n_4519), .B0 (n_2224), .Y(n_4346));
AOI21X1 g38384(.A0 (u8_mem_b3_b_127 ), .A1 (n_3879), .B0 (n_1489), .Y(n_3858));
NAND2X1 g39551(.A (n_12204), .B (u6_mem_b0_b_96 ), .Y (n_11713));
OAI21X1 g37204(.A0 (u9_rp_b1_b ), .A1 (u9_wp_b2_b ), .B0 (n_984), .Y(n_2624));
NAND2X1 g39550(.A (u7_mem_b2_b_54 ), .B (n_12650), .Y (n_4171));
NAND2X1 g37718(.A (n_4154), .B (n_3037), .Y (n_12060));
AOI21X1 g37249(.A0 (n_5359), .A1 (n_6594), .B0 (n_3958), .Y (n_5360));
AOI21X1 g37248(.A0 (n_5512), .A1 (n_6594), .B0 (n_4660), .Y (n_5513));
AOI21X1 g37247(.A0 (n_5514), .A1 (n_6594), .B0 (n_4661), .Y (n_5515));
AOI21X1 g37246(.A0 (n_5516), .A1 (n_6594), .B0 (n_4663), .Y (n_5517));
AOI21X1 g37245(.A0 (n_5518), .A1 (n_6594), .B0 (n_4664), .Y (n_5519));
MX2X1 g37244(.A (u10_mem_b1_b_148 ), .B (n_5330), .S0 (n_6475), .Y(n_5362));
AOI21X1 g37243(.A0 (n_5363), .A1 (n_6594), .B0 (n_3959), .Y (n_5364));
AOI21X1 g37242(.A0 (n_5520), .A1 (n_6594), .B0 (n_4666), .Y (n_5521));
MX2X1 g37241(.A (u9_mem_b2_b_117 ), .B (n_4764), .S0 (n_6898), .Y(n_4765));
AOI21X1 g37240(.A0 (n_5365), .A1 (n_5371), .B0 (n_3955), .Y (n_5366));
OR2X1 g41239(.A (n_697), .B (n_529), .Y (n_1484));
NOR2X1 g41238(.A (u10_rp_b2_b ), .B (u10_wp_b3_b ), .Y (n_514));
OAI21X1 g33009(.A0 (n_7264), .A1 (n_7100), .B0 (n_12609), .Y(n_9804));
OAI21X1 g33008(.A0 (n_7265), .A1 (n_7101), .B0 (n_12609), .Y(n_12835));
OAI21X1 g33005(.A0 (n_7129), .A1 (n_6996), .B0 (n_12609), .Y(n_9808));
OAI21X1 g33004(.A0 (n_7130), .A1 (n_7162), .B0 (n_12609), .Y(n_9810));
OAI21X1 g33007(.A0 (n_7127), .A1 (n_6994), .B0 (n_12609), .Y(n_9806));
OAI21X1 g33006(.A0 (n_7128), .A1 (n_7173), .B0 (n_12609), .Y(n_9807));
OAI21X1 g33001(.A0 (n_7268), .A1 (n_7102), .B0 (n_12609), .Y(n_9813));
OAI21X1 g33003(.A0 (n_7266), .A1 (n_6997), .B0 (n_12609), .Y(n_9811));
OAI21X1 g33002(.A0 (n_7132), .A1 (n_6993), .B0 (n_12609), .Y(n_9812));
NOR2X1 g45512(.A (oc0_cfg_965), .B (n_925), .Y (n_12114));
NAND2X1 g39365(.A (n_12679), .B (u5_mem_b0_b_115 ), .Y (n_3238));
NAND4X1 g45513(.A (n_12833), .B (n_12834), .C (n_3019), .D (n_1515),.Y (n_12116));
AOI21X1 g38503(.A0 (u5_mem_b2_b_33 ), .A1 (n_4370), .B0 (n_2132), .Y(n_4308));
BUFX3 g45511(.A (n_12114), .Y (n_12115));
INVX1 g41958(.A (u7_wp_b2_b ), .Y (n_1443));
INVX4 g40942(.A (n_1159), .Y (n_3911));
NAND2X1 g40943(.A (n_4738), .B (n_625), .Y (n_1159));
INVX2 g40944(.A (n_12664), .Y (n_7077));
NAND2X1 g45517(.A (n_6763), .B (u7_rp_b0_b ), .Y (n_12120));
INVX1 g41956(.A (u14_n_135), .Y (n_1119));
NOR2X1 g41092(.A (n_708), .B (u10_wp_b2_b ), .Y (n_832));
CLKBUFX1 g41091(.A (n_832), .Y (n_5407));
OAI21X1 g45515(.A0 (n_12124), .A1 (n_12125), .B0 (n_12161), .Y(n_12193));
INVX1 g41954(.A (n_8528), .Y (n_924));
NAND2X1 g41099(.A (n_8550), .B (n_503), .Y (n_9589));
INVX1 g41955(.A (u9_mem_b1_b_134 ), .Y (n_6884));
INVX1 g41952(.A (u9_mem_b2_b_93 ), .Y (n_6900));
NOR2X1 g34273(.A (u8_wp_b0_b ), .B (n_7976), .Y (n_8248));
NOR2X1 g39369(.A (n_3332), .B (n_2767), .Y (n_3234));
AOI21X1 g35469(.A0 (i3_re), .A1 (u9_rp_b1_b ), .B0 (n_6708), .Y(n_7152));
NAND3X1 g30108(.A (n_10992), .B (n_9998), .C (n_10332), .Y (n_10993));
INVX1 g41986(.A (u11_mem_b1_b_145 ), .Y (n_1599));
NAND2X1 g36991(.A (n_1569), .B (n_1832), .Y (n_4002));
NAND2X1 g34271(.A (u3_mem_b2_b_46 ), .B (n_8101), .Y (n_8129));
MX2X1 g38677(.A (u8_mem_b0_b_118 ), .B (wb_din_688), .S0 (n_3826), .Y(n_3686));
NAND2X1 g31717(.A (n_5494), .B (n_10385), .Y (n_10356));
NAND2X1 g31716(.A (n_5582), .B (n_10391), .Y (n_10357));
NAND2X1 g31715(.A (n_2538), .B (n_10065), .Y (n_9977));
NAND2X1 g31714(.A (n_5580), .B (n_10391), .Y (n_10358));
NAND2X1 g31713(.A (n_215), .B (n_10081), .Y (n_9978));
NAND2X1 g31712(.A (n_143), .B (n_10065), .Y (n_9979));
NAND2X1 g31711(.A (n_1676), .B (n_10065), .Y (n_9980));
NAND2X1 g31710(.A (n_147), .B (n_10010), .Y (n_9981));
MX2X1 g36042(.A (n_6570), .B (n_6569), .S0 (n_6594), .Y (n_6571));
INVX1 g42762(.A (u9_mem_b0_b_152 ), .Y (n_6857));
INVX1 g42763(.A (u10_mem_b3_b_83 ), .Y (n_5357));
INVX1 g42764(.A (n_836), .Y (n_4713));
NAND2X1 g31719(.A (n_196), .B (n_10010), .Y (n_9976));
AOI21X1 g35653(.A0 (n_11986), .A1 (n_11987), .B0 (n_7214), .Y(n_7215));
AOI21X1 g35650(.A0 (n_5905), .A1 (n_5747), .B0 (n_7120), .Y (n_7121));
AOI21X1 g35651(.A0 (n_6286), .A1 (n_5744), .B0 (n_7212), .Y (n_7216));
OAI21X1 g35872(.A0 (n_5565), .A1 (n_7115), .B0 (n_5887), .Y (n_6998));
AOI21X1 g35657(.A0 (n_5908), .A1 (n_5758), .B0 (n_7212), .Y (n_7118));
NAND2X1 g34270(.A (u8_mem_b3_b_129 ), .B (n_7976), .Y (n_8130));
AOI21X1 g35655(.A0 (n_6292), .A1 (n_5743), .B0 (n_7212), .Y (n_7213));
NAND4X1 g36998(.A (n_12817), .B (n_12818), .C (n_4157), .D (n_2417),.Y (n_6781));
AOI21X1 g35658(.A0 (n_6218), .A1 (n_6282), .B0 (n_7214), .Y (n_7211));
AOI21X1 g35659(.A0 (n_6166), .A1 (n_6280), .B0 (n_7214), .Y (n_7210));
OAI21X1 g35878(.A0 (n_5714), .A1 (n_7115), .B0 (n_6243), .Y (n_7173));
OAI21X1 g35879(.A0 (n_5562), .A1 (n_7115), .B0 (n_5875), .Y (n_6994));
AOI21X1 g31797(.A0 (n_5394), .A1 (n_9483), .B0 (n_9496), .Y (n_9484));
OAI21X1 g31024(.A0 (n_5336), .A1 (n_10820), .B0 (n_10388), .Y(n_10895));
MX2X1 g40426(.A (crac_din_695), .B (in_slt_834), .S0 (n_1036), .Y(n_1034));
NOR2X1 g39312(.A (n_3332), .B (n_2782), .Y (n_3285));
AOI21X1 g31795(.A0 (n_5400), .A1 (n_9546), .B0 (n_9558), .Y (n_9547));
INVX1 g42544(.A (u9_mem_b3_b_74 ), .Y (n_6089));
INVX1 g42545(.A (u10_mem_b3_b_68 ), .Y (n_6595));
AOI21X1 g31794(.A0 (n_4070), .A1 (n_9486), .B0 (n_9497), .Y (n_9487));
NAND2X1 g34277(.A (u3_mem_b2_b_52 ), .B (n_8101), .Y (n_8123));
INVX1 g42541(.A (u10_mem_b0_b_173 ), .Y (n_1685));
INVX1 g42542(.A (u11_mem_b3_b_78 ), .Y (n_5488));
INVX1 g42543(.A (u9_mem_b2_b_97 ), .Y (n_6647));
AOI21X1 g31793(.A0 (n_5396), .A1 (n_9548), .B0 (n_9559), .Y (n_9549));
INVX1 g42548(.A (u11_mem_b0_b_161 ), .Y (n_6368));
INVX1 g42549(.A (n_528), .Y (n_4711));
NAND2X1 g39212(.A (n_12389), .B (u4_mem_b0_b_110 ), .Y (n_3366));
AOI21X1 g31792(.A0 (n_5398), .A1 (n_9488), .B0 (n_9498), .Y (n_9489));
OAI21X1 g31023(.A0 (n_5406), .A1 (n_10880), .B0 (n_10389), .Y(n_10896));
NAND2X1 g39311(.A (n_12721), .B (u3_mem_b0_b_96 ), .Y (n_3287));
AOI21X1 g31790(.A0 (n_10990), .A1 (n_9876), .B0 (n_10634), .Y(n_10991));
INVX1 g42052(.A (oc3_int_set_713), .Y (n_676));
NAND2X1 g39718(.A (u4_mem_b1_b_65 ), .B (n_12265), .Y (n_12830));
NOR2X1 g39717(.A (n_3332), .B (n_2864), .Y (n_2998));
NAND2X1 g39716(.A (n_3252), .B (u7_mem_b0_b_111 ), .Y (n_2999));
NAND2X1 g39715(.A (n_12721), .B (u3_mem_b0_b_97 ), .Y (n_3000));
NAND2X1 g39714(.A (u5_mem_b2_b_56 ), .B (n_12823), .Y (n_2258));
NOR2X1 g39713(.A (n_3117), .B (n_2831), .Y (n_3001));
NAND2X1 g39712(.A (u5_mem_b1_b_70 ), .B (n_3236), .Y (n_12032));
NAND2X1 g39711(.A (u3_mem_b1_b_90 ), .B (n_3316), .Y (n_3003));
NAND2X1 g39710(.A (n_12825), .B (u3_mem_b0_b_119 ), .Y (n_3004));
NAND2X1 g36839(.A (n_1204), .B (n_2368), .Y (n_1813));
NAND4X1 g36838(.A (n_4113), .B (n_2489), .C (n_3112), .D (n_1524), .Y(n_6209));
NAND2X1 g39419(.A (u5_mem_b2_b_32 ), .B (n_12823), .Y (n_12799));
NAND2X1 g36832(.A (n_2527), .B (n_3892), .Y (n_4821));
INVX1 g36830(.A (n_6777), .Y (n_6084));
INVX1 g36835(.A (n_12354), .Y (n_6082));
NAND2X1 g34275(.A (u8_mem_b2_b_41 ), .B (n_7976), .Y (n_8125));
NOR2X1 g35454(.A (n_844), .B (n_632), .Y (n_7379));
NAND2X1 g34274(.A (u8_mem_b1_b_63 ), .B (n_7976), .Y (n_8126));
NOR2X1 g35455(.A (n_829), .B (n_631), .Y (n_7378));
NAND2X1 g39364(.A (u5_mem_b1_b_84 ), .B (n_3239), .Y (n_3240));
NOR2X1 g35456(.A (n_807), .B (n_630), .Y (n_7434));
NAND2X1 g39414(.A (in_slt_401), .B (n_3415), .Y (n_3195));
INVX1 g35457(.A (n_7385), .Y (n_865));
NAND2X1 g39415(.A (n_3255), .B (u5_mem_b0_b_93 ), .Y (n_3193));
NAND2X1 g41017(.A (u9_rp_b1_b ), .B (n_121), .Y (n_1221));
NAND2X1 g34299(.A (u3_mem_b3_b_135 ), .B (n_8101), .Y (n_8096));
NAND2X1 g34298(.A (u3_mem_b3_b_134 ), .B (n_8097), .Y (n_8098));
OAI21X1 g33829(.A0 (n_5119), .A1 (n_9034), .B0 (n_7693), .Y (n_9035));
OAI21X1 g33828(.A0 (n_4894), .A1 (n_9036), .B0 (n_7695), .Y (n_9037));
NAND2X1 g34295(.A (u3_mem_b3_b_131 ), .B (n_8101), .Y (n_8102));
NAND2X1 g34294(.A (u3_mem_b3_b ), .B (n_8101), .Y (n_8104));
NAND2X1 g34297(.A (u3_mem_b3_b_133 ), .B (n_8097), .Y (n_8099));
NAND2X1 g34296(.A (u3_mem_b3_b_132 ), .B (n_8101), .Y (n_8100));
OAI21X1 g33823(.A0 (n_4975), .A1 (n_9043), .B0 (n_7702), .Y (n_9044));
NAND2X1 g34290(.A (u3_mem_b2_b_34 ), .B (n_8101), .Y (n_8109));
NAND2X1 g34293(.A (u3_mem_b2_b_37 ), .B (n_8101), .Y (n_8105));
NAND2X1 g34292(.A (u3_mem_b2_b_36 ), .B (n_8141), .Y (n_8106));
NAND2X1 g38920(.A (u3_mem_b3_b_137 ), .B (n_1517), .Y (n_1348));
NAND2X1 g45792(.A (n_2330), .B (u7_mem_b0_b_94 ), .Y (n_12507));
NAND2X1 g34278(.A (u3_mem_b2_b_53 ), .B (n_8141), .Y (n_8122));
NOR2X1 g39511(.A (n_3117), .B (n_2792), .Y (n_3131));
OAI21X1 g33580(.A0 (n_5094), .A1 (n_9346), .B0 (n_7973), .Y (n_9347));
OAI21X1 g33581(.A0 (n_5092), .A1 (n_9346), .B0 (n_7972), .Y (n_9345));
NAND2X1 g39209(.A (n_12389), .B (u4_mem_b0_b_100 ), .Y (n_11646));
OAI21X1 g33582(.A0 (n_5091), .A1 (n_9346), .B0 (n_7971), .Y (n_9344));
NAND2X1 g39208(.A (in_slt_400), .B (n_3415), .Y (n_3373));
AOI21X1 g32990(.A0 (i4_dout_595), .A1 (n_7468), .B0 (n_8485), .Y(n_9454));
OAI21X1 g32991(.A0 (n_7326), .A1 (n_7292), .B0 (n_12149), .Y(n_11948));
OAI21X1 g32992(.A0 (n_7325), .A1 (n_7196), .B0 (n_12149), .Y(n_12012));
OAI21X1 g33583(.A0 (n_5090), .A1 (n_8318), .B0 (n_7970), .Y (n_9343));
OAI21X1 g32995(.A0 (n_7320), .A1 (n_7104), .B0 (n_9885), .Y(n_12042));
OAI21X1 g32996(.A0 (n_7319), .A1 (n_7194), .B0 (n_9885), .Y(n_11950));
OAI21X1 g32997(.A0 (n_7273), .A1 (n_7103), .B0 (n_12149), .Y(n_11980));
OAI21X1 g32999(.A0 (n_7270), .A1 (n_7201), .B0 (n_9885), .Y(n_11674));
OAI21X1 g33585(.A0 (n_5088), .A1 (n_8318), .B0 (n_7968), .Y (n_9340));
NAND2X1 g39205(.A (u4_mem_b2_b_33 ), .B (n_12087), .Y (n_3376));
OAI21X1 g33586(.A0 (n_5087), .A1 (n_8318), .B0 (n_7967), .Y (n_9339));
INVX1 g39054(.A (n_3985), .Y (n_1910));
OAI21X1 g33587(.A0 (n_5086), .A1 (n_9336), .B0 (n_7966), .Y (n_9338));
INVX1 g40780(.A (n_1172), .Y (n_2096));
NAND2X1 g39206(.A (u3_mem_b1_b_76 ), .B (n_3316), .Y (n_3375));
NAND2X1 g39512(.A (u5_mem_b1_b_85 ), .B (n_3239), .Y (n_3130));
BUFX3 g39055(.A (n_3985), .Y (n_4726));
NAND2X1 g39203(.A (n_3252), .B (u7_mem_b0_b ), .Y (n_3378));
MX2X1 g37295(.A (u11_mem_b2_b_109 ), .B (n_5315), .S0 (n_5312), .Y(n_5316));
NAND2X1 g32668(.A (n_401), .B (n_10645), .Y (n_11969));
NAND2X1 g32669(.A (n_259), .B (n_10645), .Y (n_11953));
MX2X1 g31248(.A (n_6405), .B (n_6404), .S0 (n_10308), .Y (n_10174));
NAND2X1 g32662(.A (n_166), .B (n_9931), .Y (n_12816));
NAND2X1 g32663(.A (n_266), .B (n_9931), .Y (n_9915));
NAND2X1 g32660(.A (n_262), .B (n_9931), .Y (n_12812));
NAND2X1 g32661(.A (n_234), .B (n_9931), .Y (n_12814));
NAND2X1 g32666(.A (n_387), .B (n_10645), .Y (n_11965));
NAND2X1 g32667(.A (n_229), .B (n_10645), .Y (n_11971));
NAND2X1 g32664(.A (n_264), .B (n_9931), .Y (n_9914));
NAND2X1 g32665(.A (n_9876), .B (n_1873), .Y (n_11108));
INVX1 g37012(.A (n_6814), .Y (n_6073));
NAND4X1 g37013(.A (n_11654), .B (n_11655), .C (n_1808), .D (n_11476),.Y (n_6814));
INVX1 g37010(.A (n_6167), .Y (n_5700));
NAND4X1 g37011(.A (n_3014), .B (n_3287), .C (n_2878), .D (n_1532), .Y(n_6167));
INVX1 g37016(.A (n_5823), .Y (n_5546));
NAND4X1 g37017(.A (n_11668), .B (n_11669), .C (n_2253), .D (n_2386),.Y (n_5823));
NAND4X1 g37014(.A (n_1347), .B (n_2999), .C (n_4217), .D (n_3452), .Y(n_5699));
NAND2X1 g37015(.A (n_2535), .B (n_2510), .Y (n_4807));
INVX1 g37018(.A (n_6174), .Y (n_5698));
NAND4X1 g37019(.A (n_3181), .B (n_2859), .C (n_2996), .D (n_1348), .Y(n_6174));
AND2X1 g36631(.A (n_3968), .B (n_4707), .Y (n_5590));
OAI21X1 g36630(.A0 (n_12851), .A1 (n_12852), .B0 (u4_rp_b0_b ), .Y(n_6129));
OAI21X1 g36633(.A0 (n_4609), .A1 (n_5222), .B0 (n_6134), .Y (n_6127));
OAI21X1 g36632(.A0 (n_4553), .A1 (n_5173), .B0 (n_6152), .Y (n_5790));
AOI21X1 g36635(.A0 (n_5591), .A1 (n_5788), .B0 (n_5275), .Y (n_5789));
OAI21X1 g36634(.A0 (n_4608), .A1 (n_5220), .B0 (n_6131), .Y (n_6126));
AOI21X1 g36637(.A0 (n_5591), .A1 (ic2_cfg_1049), .B0 (n_4723), .Y(n_5587));
AOI21X1 g36636(.A0 (n_5591), .A1 (n_5588), .B0 (n_4725), .Y (n_5589));
AOI21X1 g36638(.A0 (n_5591), .A1 (ic2_cfg_1050), .B0 (n_4720), .Y(n_5586));
INVX1 g42768(.A (oc5_cfg_1015), .Y (n_590));
NAND2X1 g39514(.A (n_3339), .B (in_slt_428), .Y (n_5290));
NOR2X1 g39510(.A (n_3008), .B (n_1488), .Y (n_1273));
NAND2X1 g34352(.A (u4_mem_b1_b_71 ), .B (n_7984), .Y (n_8052));
OAI22X1 g30743(.A0 (n_10950), .A1 (n_5566), .B0 (out_slt6), .B1(n_10949), .Y (n_10952));
OAI22X1 g30742(.A0 (n_10954), .A1 (n_6080), .B0 (n_10953), .B1(out_slt_84), .Y (n_10955));
OAI22X1 g30741(.A0 (n_10954), .A1 (n_6077), .B0 (out_slt4), .B1(n_10953), .Y (n_10956));
AOI21X1 g30740(.A0 (n_9695), .A1 (n_9651), .B0 (n_9586), .Y (n_9696));
OAI22X1 g30747(.A0 (n_11105), .A1 (n_5697), .B0 (out_slt8), .B1(n_11104), .Y (n_11107));
OAI22X1 g30746(.A0 (n_11109), .A1 (n_5703), .B0 (n_11108), .B1(out_slt_122), .Y (n_11110));
OAI22X1 g30745(.A0 (n_11109), .A1 (n_5556), .B0 (out_slt7), .B1(n_11108), .Y (n_11111));
OAI22X1 g30744(.A0 (n_10950), .A1 (n_5558), .B0 (n_10949), .B1(out_slt_103), .Y (n_10951));
OAI22X1 g30749(.A0 (n_11100), .A1 (n_5686), .B0 (out_slt3), .B1(n_11099), .Y (n_11103));
OAI22X1 g30748(.A0 (n_11105), .A1 (n_5715), .B0 (n_11104), .B1(out_slt_141), .Y (n_11106));
NAND2X1 g39517(.A (u3_mem_b2_b_29 ), .B (n_12619), .Y (n_3126));
MX2X1 g38598(.A (u8_mem_b0_b_101 ), .B (wb_din_671), .S0 (n_3826), .Y(n_3814));
MX2X1 g38599(.A (u3_mem_b0_b_104 ), .B (wb_din_674), .S0 (n_3807), .Y(n_3813));
MX2X1 g38596(.A (u8_mem_b0_b_102 ), .B (wb_din_672), .S0 (n_3826), .Y(n_3817));
MX2X1 g38597(.A (u3_mem_b0_b_107 ), .B (wb_din_677), .S0 (n_3807), .Y(n_3815));
MX2X1 g38594(.A (u3_mem_b0_b_92 ), .B (wb_din_662), .S0 (n_858), .Y(n_3820));
MX2X1 g38595(.A (u8_mem_b0_b_103 ), .B (wb_din_673), .S0 (n_3826), .Y(n_3818));
MX2X1 g38592(.A (u3_mem_b0_b_109 ), .B (wb_din_679), .S0 (n_3807), .Y(n_3823));
MX2X1 g38593(.A (u8_mem_b0_b_121 ), .B (wb_din_691), .S0 (n_3826), .Y(n_3822));
MX2X1 g38590(.A (u8_mem_b0_b_107 ), .B (wb_din_677), .S0 (n_3826), .Y(n_3825));
MX2X1 g38591(.A (u8_mem_b0_b_105 ), .B (wb_din_675), .S0 (n_3826), .Y(n_3824));
NOR2X1 g39516(.A (n_4996), .B (n_2790), .Y (n_3128));
NOR2X1 g39682(.A (n_3117), .B (n_2801), .Y (n_3023));
INVX4 g40867(.A (n_1019), .Y (n_2477));
OR2X1 g35458(.A (n_632), .B (n_11563), .Y (n_7385));
NAND2X1 g39684(.A (u4_mem_b1_b_77 ), .B (n_12250), .Y (n_4144));
INVX2 g39052(.A (n_1910), .Y (n_3979));
NOR2X1 g41394(.A (n_12332), .B (n_12330), .Y (n_846));
INVX1 g41396(.A (n_9717), .Y (n_7120));
NAND2X1 g41390(.A (u10_wp_b1_b ), .B (u10_wp_b2_b ), .Y (n_1067));
BUFX3 g41391(.A (n_846), .Y (n_1538));
INVX1 g41392(.A (n_1546), .Y (n_1068));
BUFX3 g41393(.A (n_846), .Y (n_1546));
INVX1 g35459(.A (n_7382), .Y (n_864));
INVX1 g41399(.A (n_9717), .Y (n_7212));
NAND2X1 g38926(.A (u7_mem_b3_b_133 ), .B (n_1538), .Y (n_1530));
MX2X1 g31266(.A (n_5474), .B (n_2500), .S0 (n_10267), .Y (n_10154));
MX2X1 g31368(.A (u10_din_tmp_48), .B (in_slt_429), .S0 (n_9860), .Y(n_9865));
MX2X1 g31369(.A (u10_din_tmp_49), .B (in_slt_430), .S0 (n_9860), .Y(n_9863));
MX2X1 g31366(.A (u9_din_tmp_50), .B (in_slt_409), .S0 (n_9777), .Y(n_9770));
MX2X1 g31367(.A (u10_din_tmp_47), .B (in_slt_428), .S0 (n_9860), .Y(n_9867));
MX2X1 g31364(.A (u9_din_tmp_48), .B (in_slt_407), .S0 (n_9777), .Y(n_9772));
MX2X1 g31365(.A (u9_din_tmp_49), .B (in_slt_408), .S0 (n_9777), .Y(n_9771));
MX2X1 g31362(.A (u9_din_tmp_46), .B (in_slt_405), .S0 (n_9777), .Y(n_9774));
MX2X1 g31363(.A (u9_din_tmp_47), .B (in_slt_406), .S0 (n_9777), .Y(n_9773));
MX2X1 g31360(.A (u9_din_tmp_44), .B (in_slt_403), .S0 (n_9777), .Y(n_9776));
MX2X1 g31361(.A (u9_din_tmp_45), .B (in_slt_404), .S0 (n_9777), .Y(n_9775));
AOI22X1 g37900(.A0 (n_2344), .A1 (in_slt_437), .B0 (n_2302), .B1(in_slt_425), .Y (n_5422));
AOI22X1 g37901(.A0 (u11_din_tmp_42), .A1 (n_4560), .B0 (n_4097), .B1(in_slt_443), .Y (n_3898));
AOI22X1 g37902(.A0 (u10_din_tmp_42), .A1 (n_2302), .B0 (n_3911), .B1(in_slt_421), .Y (n_2511));
NAND2X1 g37903(.A (n_3557), .B (n_3013), .Y (n_4569));
AOI22X1 g37904(.A0 (n_2558), .A1 (n_6384), .B0 (n_6468), .B1(n_1839), .Y (n_1840));
AOI22X1 g37905(.A0 (n_6476), .A1 (n_940), .B0 (n_6601), .B1 (n_1316),.Y (n_2510));
AOI22X1 g37906(.A0 (u11_din_tmp_43), .A1 (n_4560), .B0 (n_4097), .B1(in_slt_444), .Y (n_3896));
NAND2X1 g37907(.A (n_3530), .B (n_3109), .Y (n_4568));
AOI22X1 g37908(.A0 (u11_din_tmp_44), .A1 (n_4560), .B0 (n_4097), .B1(in_slt_445), .Y (n_3895));
AOI22X1 g37909(.A0 (n_2502), .A1 (n_1562), .B0 (n_1561), .B1(n_1835), .Y (n_1563));
INVX1 g39513(.A (n_5290), .Y (n_4178));
MX2X1 g33210(.A (u13_intm_r_b28_b ), .B (wb_din_688), .S0 (n_8519), .Y(n_8496));
MX2X1 g33211(.A (u13_intm_r_b2_b ), .B (wb_din_662), .S0 (n_8519), .Y(n_8494));
MX2X1 g33212(.A (u13_intm_r_b3_b ), .B (wb_din_663), .S0 (n_8519), .Y(n_8493));
MX2X1 g33213(.A (u13_intm_r_b4_b ), .B (wb_din_664), .S0 (n_8519), .Y(n_8492));
MX2X1 g33214(.A (u13_intm_r_b5_b ), .B (wb_din_665), .S0 (n_8519), .Y(n_8491));
MX2X1 g33215(.A (u13_intm_r_b6_b ), .B (wb_din_666), .S0 (n_8519), .Y(n_8490));
MX2X1 g33216(.A (u13_intm_r_b7_b ), .B (wb_din_667), .S0 (n_8519), .Y(n_8489));
MX2X1 g33217(.A (u13_intm_r_b8_b ), .B (wb_din_668), .S0 (n_8519), .Y(n_8488));
MX2X1 g33218(.A (u13_intm_r_b9_b ), .B (wb_din_669), .S0 (n_8519), .Y(n_8487));
NOR2X1 g41179(.A (n_4710), .B (n_836), .Y (n_1049));
NAND2X1 g34848(.A (u8_mem_b1_b_68 ), .B (n_7976), .Y (n_7586));
NAND2X1 g34849(.A (u3_mem_b1_b_75 ), .B (n_8141), .Y (n_7585));
INVX1 g42159(.A (u10_mem_b1_b_129 ), .Y (n_6468));
INVX1 g42158(.A (u11_mem_b1_b_149 ), .Y (n_1580));
NAND2X1 g34840(.A (u8_mem_b1_b_89 ), .B (n_7976), .Y (n_7594));
NAND2X1 g34841(.A (u3_mem_b1_b_71 ), .B (n_8101), .Y (n_7593));
NAND2X1 g34842(.A (u8_mem_b1_b_90 ), .B (n_7976), .Y (n_7592));
NAND2X1 g34843(.A (u3_mem_b1_b_72 ), .B (n_8101), .Y (n_7591));
NAND2X1 g34844(.A (u8_mem_b1_b_64 ), .B (n_7976), .Y (n_7590));
NAND2X1 g34845(.A (u3_mem_b1_b_73 ), .B (n_8141), .Y (n_7589));
NAND2X1 g34846(.A (u8_mem_b1_b_65 ), .B (n_7976), .Y (n_7588));
NAND2X1 g34847(.A (u8_mem_b1_b_67 ), .B (n_7976), .Y (n_7587));
NAND2X1 g39942(.A (n_11789), .B (u8_mem_b0_b_95 ), .Y (n_2861));
NAND2X1 g39943(.A (n_3259), .B (u5_mem_b0_b_107 ), .Y (n_12857));
NAND2X1 g39940(.A (n_3259), .B (u5_mem_b0_b_105 ), .Y (n_12841));
NAND2X1 g39941(.A (n_2491), .B (u7_mem_b0_b_99 ), .Y (n_2493));
NOR2X1 g39946(.A (n_3089), .B (n_2716), .Y (n_2858));
NAND2X1 g39947(.A (u5_mem_b1_b_89 ), .B (n_3236), .Y (n_2857));
NAND2X1 g39944(.A (n_12721), .B (u3_mem_b0_b_106 ), .Y (n_2859));
NAND2X2 g39945(.A (n_1367), .B (u8_rp_b3_b ), .Y (n_4829));
NAND2X1 g39948(.A (u5_mem_b2_b_58 ), .B (n_12823), .Y (n_2231));
NAND2X1 g39949(.A (n_12825), .B (u3_mem_b0_b_116 ), .Y (n_2856));
INVX1 g45862(.A (oc5_cfg), .Y (n_12584));
OAI21X1 g33456(.A0 (n_4522), .A1 (n_8097), .B0 (n_8121), .Y (n_8404));
OAI21X1 g33457(.A0 (n_4341), .A1 (n_8856), .B0 (n_8120), .Y (n_8403));
OAI21X1 g33454(.A0 (n_4524), .A1 (n_8911), .B0 (n_8060), .Y (n_8406));
NAND2X1 g39366(.A (u5_mem_b1_b_72 ), .B (n_3236), .Y (n_12798));
NAND2X1 g39367(.A (u7_mem_b1_b ), .B (n_4130), .Y (n_4199));
OAI21X1 g33771(.A0 (n_4988), .A1 (n_9110), .B0 (n_7756), .Y (n_9108));
OAI21X1 g33455(.A0 (n_4320), .A1 (n_8101), .B0 (n_8123), .Y (n_8405));
NOR2X1 g39362(.A (n_4961), .B (n_2818), .Y (n_3242));
NAND2X1 g39363(.A (u5_mem_b2_b_53 ), .B (n_12823), .Y (n_2317));
NAND2X1 g39360(.A (n_3259), .B (u5_mem_b0_b_102 ), .Y (n_12853));
NAND2X1 g39361(.A (u5_mem_b2_b_40 ), .B (n_12823), .Y (n_12854));
NAND2X1 g34332(.A (u8_mem_b2_b_34 ), .B (n_7976), .Y (n_8070));
NAND2X1 g45925(.A (n_12666), .B (n_12667), .Y (n_12668));
NOR2X1 g39368(.A (n_3332), .B (n_3008), .Y (n_3235));
OAI21X1 g33453(.A0 (n_4474), .A1 (n_8393), .B0 (n_7946), .Y (n_8407));
OR2X1 g30109(.A (u13_ints_r_b20_b ), .B (ic0_int_set), .Y (n_9693));
AOI21X1 g35468(.A0 (i4_dout_613), .A1 (n_7468), .B0 (n_7138), .Y(n_7336));
NAND4X1 g36997(.A (n_4158), .B (n_3125), .C (n_2274), .D (n_2407), .Y(n_5829));
OAI21X1 g33450(.A0 (n_4347), .A1 (n_8911), .B0 (n_8127), .Y (n_8411));
INVX1 g36992(.A (n_5847), .Y (n_5549));
NAND4X1 g36993(.A (n_11703), .B (n_11704), .C (n_2264), .D (n_2423),.Y (n_5847));
MX2X1 g40421(.A (crac_din_696), .B (in_slt_835), .S0 (n_1036), .Y(n_1197));
OR2X1 g35460(.A (n_11597), .B (n_631), .Y (n_7382));
MX2X1 g34014(.A (u5_mem_b0_b ), .B (n_3741), .S0 (n_7496), .Y(n_8809));
NAND2X1 g34331(.A (n_6703), .B (n_7460), .Y (n_8237));
AOI21X1 g35465(.A0 (u11_rp_b1_b ), .A1 (i6_re), .B0 (n_6750), .Y(n_7153));
NAND3X1 g35464(.A (n_6061), .B (n_729), .C (n_730), .Y (n_7021));
AOI21X1 g35467(.A0 (i4_dout_612), .A1 (n_7468), .B0 (n_7139), .Y(n_7337));
NOR2X1 g35466(.A (n_6043), .B (n_7019), .Y (n_7020));
NAND2X1 g34592(.A (u3_mem_b2_b_48 ), .B (n_8141), .Y (n_7835));
NAND2X1 g34593(.A (u3_mem_b3_b_130 ), .B (n_8101), .Y (n_7834));
NAND2X1 g34590(.A (u8_mem_b3_b_127 ), .B (n_7976), .Y (n_7837));
NAND2X1 g34591(.A (u8_mem_b3_b_130 ), .B (n_7976), .Y (n_7836));
NOR2X1 g34596(.A (o4_status_972), .B (n_458), .Y (n_9548));
NOR2X1 g34597(.A (o6_status_982), .B (n_447), .Y (n_9486));
NAND2X1 g34594(.A (u8_mem_b3_b_128 ), .B (n_7976), .Y (n_7833));
NOR2X1 g34595(.A (o3_status_962), .B (n_459), .Y (n_9488));
NAND2X1 g34598(.A (u6_mem_b1_b ), .B (n_7758), .Y (n_7832));
NAND2X1 g34599(.A (u6_mem_b1_b_69 ), .B (n_7758), .Y (n_7831));
INVX8 g32857(.A (n_9726), .Y (n_10137));
OAI21X1 g33458(.A0 (n_4521), .A1 (n_8101), .B0 (n_8119), .Y (n_8402));
OAI21X1 g33459(.A0 (n_4520), .A1 (n_8440), .B0 (n_8117), .Y (n_8401));
NAND2X1 g31642(.A (n_5352), .B (n_10010), .Y (n_10002));
NAND2X1 g40698(.A (n_4703), .B (n_872), .Y (n_7526));
NAND2X1 g45810(.A (n_12530), .B (n_12531), .Y (n_12532));
NAND2X1 g34336(.A (u8_mem_b2_b_32 ), .B (n_7976), .Y (n_8067));
NAND2X1 g34337(.A (u3_mem_b2_b_51 ), .B (n_8101), .Y (n_8066));
NAND2X1 g34334(.A (u3_mem_b1_b_68 ), .B (n_8101), .Y (n_8069));
NAND2X1 g34335(.A (u3_mem_b1_b_87 ), .B (n_8101), .Y (n_8068));
OAI21X1 g33452(.A0 (n_5156), .A1 (n_8911), .B0 (n_8167), .Y (n_8408));
NAND2X1 g34333(.A (n_6702), .B (n_7471), .Y (n_8236));
NAND2X1 g34330(.A (u8_mem_b2_b_36 ), .B (n_7976), .Y (n_8072));
OAI21X1 g33451(.A0 (n_4526), .A1 (n_8097), .B0 (n_7724), .Y (n_8410));
NAND2X1 g34338(.A (u3_mem_b3_b_126 ), .B (n_8141), .Y (n_8065));
NAND2X1 g34339(.A (u3_mem_b1_b_67 ), .B (n_8141), .Y (n_8064));

endmodule